`timescale 1ns / 1ns

module Mac(
  input          clock,
  input          reset,
  input  [399:0] io_a,
  input  [399:0] io_b,
  input          io_rdy,
  output [31:0]  io_q,
  output         io_v
);
  wire [15:0] a_0;
  wire [15:0] b_0;
  wire [15:0] a_1;
  wire [15:0] b_1;
  wire [15:0] a_2;
  wire [15:0] b_2;
  wire [15:0] a_3;
  wire [15:0] b_3;
  wire [15:0] a_4;
  wire [15:0] b_4;
  wire [15:0] a_5;
  wire [15:0] b_5;
  wire [15:0] a_6;
  wire [15:0] b_6;
  wire [15:0] a_7;
  wire [15:0] b_7;
  wire [15:0] a_8;
  wire [15:0] b_8;
  wire [15:0] a_9;
  wire [15:0] b_9;
  wire [15:0] a_10;
  wire [15:0] b_10;
  wire [15:0] a_11;
  wire [15:0] b_11;
  wire [15:0] a_12;
  wire [15:0] b_12;
  wire [15:0] a_13;
  wire [15:0] b_13;
  wire [15:0] a_14;
  wire [15:0] b_14;
  wire [15:0] a_15;
  wire [15:0] b_15;
  wire [15:0] a_16;
  wire [15:0] b_16;
  wire [15:0] a_17;
  wire [15:0] b_17;
  wire [15:0] a_18;
  wire [15:0] b_18;
  wire [15:0] a_19;
  wire [15:0] b_19;
  wire [15:0] a_20;
  wire [15:0] b_20;
  wire [15:0] a_21;
  wire [15:0] b_21;
  wire [15:0] a_22;
  wire [15:0] b_22;
  wire [15:0] a_23;
  wire [15:0] b_23;
  wire [15:0] a_24;
  wire [15:0] b_24;
  reg [31:0] sum;
  reg [31:0] _RAND_0;
  reg [4:0] i;
  reg [31:0] _RAND_1;
  wire  _T_53;
  wire  _T_54;
  wire [15:0] _GEN_1;
  wire [15:0] _GEN_2;
  wire [15:0] _GEN_3;
  wire [15:0] _GEN_4;
  wire [15:0] _GEN_5;
  wire [15:0] _GEN_6;
  wire [15:0] _GEN_7;
  wire [15:0] _GEN_8;
  wire [15:0] _GEN_9;
  wire [15:0] _GEN_10;
  wire [15:0] _GEN_11;
  wire [15:0] _GEN_12;
  wire [15:0] _GEN_13;
  wire [15:0] _GEN_14;
  wire [15:0] _GEN_15;
  wire [15:0] _GEN_16;
  wire [15:0] _GEN_17;
  wire [15:0] _GEN_18;
  wire [15:0] _GEN_19;
  wire [15:0] _GEN_20;
  wire [15:0] _GEN_21;
  wire [15:0] _GEN_22;
  wire [15:0] _GEN_23;
  wire [15:0] _GEN_24;
  wire [15:0] _GEN_26;
  wire [15:0] _GEN_27;
  wire [15:0] _GEN_28;
  wire [15:0] _GEN_29;
  wire [15:0] _GEN_30;
  wire [15:0] _GEN_31;
  wire [15:0] _GEN_32;
  wire [15:0] _GEN_33;
  wire [15:0] _GEN_34;
  wire [15:0] _GEN_35;
  wire [15:0] _GEN_36;
  wire [15:0] _GEN_37;
  wire [15:0] _GEN_38;
  wire [15:0] _GEN_39;
  wire [15:0] _GEN_40;
  wire [15:0] _GEN_41;
  wire [15:0] _GEN_42;
  wire [15:0] _GEN_43;
  wire [15:0] _GEN_44;
  wire [15:0] _GEN_45;
  wire [15:0] _GEN_46;
  wire [15:0] _GEN_47;
  wire [15:0] _GEN_48;
  wire [15:0] _GEN_49;
  wire [31:0] _T_50;
  wire [32:0] _T_51;
  wire [5:0] _T_52;
  wire [5:0] _GEN_50;
  wire [32:0] _GEN_51;
  wire [5:0] _GEN_52;
  wire [31:0] _GEN_54;
  wire [32:0] _GEN_55;
  wire [32:0] _GEN_56;
  wire [5:0] _GEN_57;
  assign a_0 = io_a[15:0];
  assign b_0 = io_b[15:0];
  assign a_1 = io_a[31:16];
  assign b_1 = io_b[31:16];
  assign a_2 = io_a[47:32];
  assign b_2 = io_b[47:32];
  assign a_3 = io_a[63:48];
  assign b_3 = io_b[63:48];
  assign a_4 = io_a[79:64];
  assign b_4 = io_b[79:64];
  assign a_5 = io_a[95:80];
  assign b_5 = io_b[95:80];
  assign a_6 = io_a[111:96];
  assign b_6 = io_b[111:96];
  assign a_7 = io_a[127:112];
  assign b_7 = io_b[127:112];
  assign a_8 = io_a[143:128];
  assign b_8 = io_b[143:128];
  assign a_9 = io_a[159:144];
  assign b_9 = io_b[159:144];
  assign a_10 = io_a[175:160];
  assign b_10 = io_b[175:160];
  assign a_11 = io_a[191:176];
  assign b_11 = io_b[191:176];
  assign a_12 = io_a[207:192];
  assign b_12 = io_b[207:192];
  assign a_13 = io_a[223:208];
  assign b_13 = io_b[223:208];
  assign a_14 = io_a[239:224];
  assign b_14 = io_b[239:224];
  assign a_15 = io_a[255:240];
  assign b_15 = io_b[255:240];
  assign a_16 = io_a[271:256];
  assign b_16 = io_b[271:256];
  assign a_17 = io_a[287:272];
  assign b_17 = io_b[287:272];
  assign a_18 = io_a[303:288];
  assign b_18 = io_b[303:288];
  assign a_19 = io_a[319:304];
  assign b_19 = io_b[319:304];
  assign a_20 = io_a[335:320];
  assign b_20 = io_b[335:320];
  assign a_21 = io_a[351:336];
  assign b_21 = io_b[351:336];
  assign a_22 = io_a[367:352];
  assign b_22 = io_b[367:352];
  assign a_23 = io_a[383:368];
  assign b_23 = io_b[383:368];
  assign a_24 = io_a[399:384];
  assign b_24 = io_b[399:384];
  assign _T_53 = i == 5'h19;
  assign _T_54 = i != 5'h0;
  assign _GEN_1 = 5'h1 == i ? a_1 : a_0;
  assign _GEN_2 = 5'h2 == i ? a_2 : _GEN_1;
  assign _GEN_3 = 5'h3 == i ? a_3 : _GEN_2;
  assign _GEN_4 = 5'h4 == i ? a_4 : _GEN_3;
  assign _GEN_5 = 5'h5 == i ? a_5 : _GEN_4;
  assign _GEN_6 = 5'h6 == i ? a_6 : _GEN_5;
  assign _GEN_7 = 5'h7 == i ? a_7 : _GEN_6;
  assign _GEN_8 = 5'h8 == i ? a_8 : _GEN_7;
  assign _GEN_9 = 5'h9 == i ? a_9 : _GEN_8;
  assign _GEN_10 = 5'ha == i ? a_10 : _GEN_9;
  assign _GEN_11 = 5'hb == i ? a_11 : _GEN_10;
  assign _GEN_12 = 5'hc == i ? a_12 : _GEN_11;
  assign _GEN_13 = 5'hd == i ? a_13 : _GEN_12;
  assign _GEN_14 = 5'he == i ? a_14 : _GEN_13;
  assign _GEN_15 = 5'hf == i ? a_15 : _GEN_14;
  assign _GEN_16 = 5'h10 == i ? a_16 : _GEN_15;
  assign _GEN_17 = 5'h11 == i ? a_17 : _GEN_16;
  assign _GEN_18 = 5'h12 == i ? a_18 : _GEN_17;
  assign _GEN_19 = 5'h13 == i ? a_19 : _GEN_18;
  assign _GEN_20 = 5'h14 == i ? a_20 : _GEN_19;
  assign _GEN_21 = 5'h15 == i ? a_21 : _GEN_20;
  assign _GEN_22 = 5'h16 == i ? a_22 : _GEN_21;
  assign _GEN_23 = 5'h17 == i ? a_23 : _GEN_22;
  assign _GEN_24 = 5'h18 == i ? a_24 : _GEN_23;
  assign _GEN_26 = 5'h1 == i ? b_1 : b_0;
  assign _GEN_27 = 5'h2 == i ? b_2 : _GEN_26;
  assign _GEN_28 = 5'h3 == i ? b_3 : _GEN_27;
  assign _GEN_29 = 5'h4 == i ? b_4 : _GEN_28;
  assign _GEN_30 = 5'h5 == i ? b_5 : _GEN_29;
  assign _GEN_31 = 5'h6 == i ? b_6 : _GEN_30;
  assign _GEN_32 = 5'h7 == i ? b_7 : _GEN_31;
  assign _GEN_33 = 5'h8 == i ? b_8 : _GEN_32;
  assign _GEN_34 = 5'h9 == i ? b_9 : _GEN_33;
  assign _GEN_35 = 5'ha == i ? b_10 : _GEN_34;
  assign _GEN_36 = 5'hb == i ? b_11 : _GEN_35;
  assign _GEN_37 = 5'hc == i ? b_12 : _GEN_36;
  assign _GEN_38 = 5'hd == i ? b_13 : _GEN_37;
  assign _GEN_39 = 5'he == i ? b_14 : _GEN_38;
  assign _GEN_40 = 5'hf == i ? b_15 : _GEN_39;
  assign _GEN_41 = 5'h10 == i ? b_16 : _GEN_40;
  assign _GEN_42 = 5'h11 == i ? b_17 : _GEN_41;
  assign _GEN_43 = 5'h12 == i ? b_18 : _GEN_42;
  assign _GEN_44 = 5'h13 == i ? b_19 : _GEN_43;
  assign _GEN_45 = 5'h14 == i ? b_20 : _GEN_44;
  assign _GEN_46 = 5'h15 == i ? b_21 : _GEN_45;
  assign _GEN_47 = 5'h16 == i ? b_22 : _GEN_46;
  assign _GEN_48 = 5'h17 == i ? b_23 : _GEN_47;
  assign _GEN_49 = 5'h18 == i ? b_24 : _GEN_48;
  assign _T_50 = _GEN_24 * _GEN_49;
  assign _T_51 = sum + _T_50;
  assign _T_52 = i + 5'h1;
  assign _GEN_50 = _T_54 ? _T_52 : 6'h0;
  assign _GEN_51 = _T_54 ? _T_51 : 33'h0;
  assign _GEN_52 = _T_53 ? 6'h0 : _GEN_50;
  assign _GEN_54 = _T_53 ? sum : 32'h0;
  assign _GEN_55 = _T_53 ? 33'h0 : _GEN_51;
  assign _GEN_56 = io_rdy ? _T_51 : _GEN_55;
  assign _GEN_57 = io_rdy ? _T_52 : _GEN_52;
  assign io_q = io_rdy ? 32'h0 : _GEN_54;
  assign io_v = io_rdy ? 1'h0 : _T_53;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sum = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  i = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      sum <= 32'h0;
    end else begin
      sum <= _GEN_56[31:0];
    end
    if (reset) begin
      i <= 5'h0;
    end else begin
      i <= _GEN_57[4:0];
    end
  end
endmodule
module ReLU(
  input  [31:0] io_q,
  input  [15:0] io_bias,
  input         io_v_in,
  output [15:0] io_d,
  output        io_v_out
);
  wire [15:0] qc;
  wire [16:0] _T_2;
  wire  _T_3;
  wire [16:0] _T_1;
  wire [16:0] _GEN_0;
  assign qc = io_q[15:0];
  assign _T_2 = qc + io_bias;
  assign _T_3 = _T_2 > 17'h0;
  assign _T_1 = _T_3 ? _T_2 : 17'h0;
  assign _GEN_0 = io_v_in ? _T_1 : 17'h0;
  assign io_d = _GEN_0[15:0];
  assign io_v_out = io_v_in;
endmodule
module Node(
  input          clock,
  input          reset,
  input  [399:0] io_d_in,
  input  [399:0] io_w,
  input          io_rdy,
  input  [15:0]  io_bias,
  output [15:0]  io_d_out,
  output         io_v
);
  wire  muladdc_clock;
  wire  muladdc_reset;
  wire [399:0] muladdc_io_a;
  wire [399:0] muladdc_io_b;
  wire  muladdc_io_rdy;
  wire [31:0] muladdc_io_q;
  wire  muladdc_io_v;
  wire [31:0] act_io_q;
  wire [15:0] act_io_bias;
  wire  act_io_v_in;
  wire [15:0] act_io_d;
  wire  act_io_v_out;
  Mac muladdc (
    .clock(muladdc_clock),
    .reset(muladdc_reset),
    .io_a(muladdc_io_a),
    .io_b(muladdc_io_b),
    .io_rdy(muladdc_io_rdy),
    .io_q(muladdc_io_q),
    .io_v(muladdc_io_v)
  );
  ReLU act (
    .io_q(act_io_q),
    .io_bias(act_io_bias),
    .io_v_in(act_io_v_in),
    .io_d(act_io_d),
    .io_v_out(act_io_v_out)
  );
  assign io_d_out = act_io_d;
  assign io_v = act_io_v_out;
  assign muladdc_clock = clock;
  assign muladdc_reset = reset;
  assign muladdc_io_a = io_d_in;
  assign muladdc_io_b = io_w;
  assign muladdc_io_rdy = io_rdy;
  assign act_io_q = muladdc_io_q;
  assign act_io_bias = io_bias;
  assign act_io_v_in = muladdc_io_v;
endmodule
module ConvC1(
  input          clock,
  input          reset,
  input  [399:0] io_d_in,
  input  [399:0] io_w_in_0,
  input  [399:0] io_w_in_1,
  input  [399:0] io_w_in_2,
  input  [399:0] io_w_in_3,
  input  [399:0] io_w_in_4,
  input  [399:0] io_w_in_5,
  input  [95:0]  io_bias,
  input          io_rdy,
  output [15:0]  io_d_out_0,
  output [15:0]  io_d_out_1,
  output [15:0]  io_d_out_2,
  output [15:0]  io_d_out_3,
  output [15:0]  io_d_out_4,
  output [15:0]  io_d_out_5,
  output         io_v
);
  wire  _T_clock;
  wire  _T_reset;
  wire [399:0] _T_io_d_in;
  wire [399:0] _T_io_w;
  wire  _T_io_rdy;
  wire [15:0] _T_io_bias;
  wire [15:0] _T_io_d_out;
  wire  _T_io_v;
  wire  _T_1_clock;
  wire  _T_1_reset;
  wire [399:0] _T_1_io_d_in;
  wire [399:0] _T_1_io_w;
  wire  _T_1_io_rdy;
  wire [15:0] _T_1_io_bias;
  wire [15:0] _T_1_io_d_out;
  wire  _T_1_io_v;
  wire  _T_2_clock;
  wire  _T_2_reset;
  wire [399:0] _T_2_io_d_in;
  wire [399:0] _T_2_io_w;
  wire  _T_2_io_rdy;
  wire [15:0] _T_2_io_bias;
  wire [15:0] _T_2_io_d_out;
  wire  _T_2_io_v;
  wire  _T_3_clock;
  wire  _T_3_reset;
  wire [399:0] _T_3_io_d_in;
  wire [399:0] _T_3_io_w;
  wire  _T_3_io_rdy;
  wire [15:0] _T_3_io_bias;
  wire [15:0] _T_3_io_d_out;
  wire  _T_3_io_v;
  wire  _T_4_clock;
  wire  _T_4_reset;
  wire [399:0] _T_4_io_d_in;
  wire [399:0] _T_4_io_w;
  wire  _T_4_io_rdy;
  wire [15:0] _T_4_io_bias;
  wire [15:0] _T_4_io_d_out;
  wire  _T_4_io_v;
  wire  _T_5_clock;
  wire  _T_5_reset;
  wire [399:0] _T_5_io_d_in;
  wire [399:0] _T_5_io_w;
  wire  _T_5_io_rdy;
  wire [15:0] _T_5_io_bias;
  wire [15:0] _T_5_io_d_out;
  wire  _T_5_io_v;
  wire  _T_6;
  wire  _T_7;
  wire  _T_8;
  wire  _T_9;
  Node _T (
    .clock(_T_clock),
    .reset(_T_reset),
    .io_d_in(_T_io_d_in),
    .io_w(_T_io_w),
    .io_rdy(_T_io_rdy),
    .io_bias(_T_io_bias),
    .io_d_out(_T_io_d_out),
    .io_v(_T_io_v)
  );
  Node _T_1 (
    .clock(_T_1_clock),
    .reset(_T_1_reset),
    .io_d_in(_T_1_io_d_in),
    .io_w(_T_1_io_w),
    .io_rdy(_T_1_io_rdy),
    .io_bias(_T_1_io_bias),
    .io_d_out(_T_1_io_d_out),
    .io_v(_T_1_io_v)
  );
  Node _T_2 (
    .clock(_T_2_clock),
    .reset(_T_2_reset),
    .io_d_in(_T_2_io_d_in),
    .io_w(_T_2_io_w),
    .io_rdy(_T_2_io_rdy),
    .io_bias(_T_2_io_bias),
    .io_d_out(_T_2_io_d_out),
    .io_v(_T_2_io_v)
  );
  Node _T_3 (
    .clock(_T_3_clock),
    .reset(_T_3_reset),
    .io_d_in(_T_3_io_d_in),
    .io_w(_T_3_io_w),
    .io_rdy(_T_3_io_rdy),
    .io_bias(_T_3_io_bias),
    .io_d_out(_T_3_io_d_out),
    .io_v(_T_3_io_v)
  );
  Node _T_4 (
    .clock(_T_4_clock),
    .reset(_T_4_reset),
    .io_d_in(_T_4_io_d_in),
    .io_w(_T_4_io_w),
    .io_rdy(_T_4_io_rdy),
    .io_bias(_T_4_io_bias),
    .io_d_out(_T_4_io_d_out),
    .io_v(_T_4_io_v)
  );
  Node _T_5 (
    .clock(_T_5_clock),
    .reset(_T_5_reset),
    .io_d_in(_T_5_io_d_in),
    .io_w(_T_5_io_w),
    .io_rdy(_T_5_io_rdy),
    .io_bias(_T_5_io_bias),
    .io_d_out(_T_5_io_d_out),
    .io_v(_T_5_io_v)
  );
  assign _T_6 = _T_io_v & _T_1_io_v;
  assign _T_7 = _T_6 & _T_2_io_v;
  assign _T_8 = _T_7 & _T_3_io_v;
  assign _T_9 = _T_8 & _T_4_io_v;
  assign io_d_out_0 = _T_io_d_out;
  assign io_d_out_1 = _T_1_io_d_out;
  assign io_d_out_2 = _T_2_io_d_out;
  assign io_d_out_3 = _T_3_io_d_out;
  assign io_d_out_4 = _T_4_io_d_out;
  assign io_d_out_5 = _T_5_io_d_out;
  assign io_v = _T_9 & _T_5_io_v;
  assign _T_clock = clock;
  assign _T_reset = reset;
  assign _T_io_d_in = io_d_in;
  assign _T_io_w = io_w_in_0;
  assign _T_io_rdy = io_rdy;
  assign _T_io_bias = io_bias[15:0];
  assign _T_1_clock = clock;
  assign _T_1_reset = reset;
  assign _T_1_io_d_in = io_d_in;
  assign _T_1_io_w = io_w_in_1;
  assign _T_1_io_rdy = io_rdy;
  assign _T_1_io_bias = io_bias[15:0];
  assign _T_2_clock = clock;
  assign _T_2_reset = reset;
  assign _T_2_io_d_in = io_d_in;
  assign _T_2_io_w = io_w_in_2;
  assign _T_2_io_rdy = io_rdy;
  assign _T_2_io_bias = io_bias[15:0];
  assign _T_3_clock = clock;
  assign _T_3_reset = reset;
  assign _T_3_io_d_in = io_d_in;
  assign _T_3_io_w = io_w_in_3;
  assign _T_3_io_rdy = io_rdy;
  assign _T_3_io_bias = io_bias[15:0];
  assign _T_4_clock = clock;
  assign _T_4_reset = reset;
  assign _T_4_io_d_in = io_d_in;
  assign _T_4_io_w = io_w_in_4;
  assign _T_4_io_rdy = io_rdy;
  assign _T_4_io_bias = io_bias[15:0];
  assign _T_5_clock = clock;
  assign _T_5_reset = reset;
  assign _T_5_io_d_in = io_d_in;
  assign _T_5_io_w = io_w_in_5;
  assign _T_5_io_rdy = io_rdy;
  assign _T_5_io_bias = io_bias[15:0];
endmodule
module MaxPool(
  input  [63:0] io_d_in,
  input         io_rdy,
  output [15:0] io_q,
  output        io_v
);
  wire [15:0] _T_1;
  wire [15:0] _T_2;
  wire [15:0] _T_3;
  wire [15:0] _T_4;
  wire  _T_5;
  wire [15:0] _GEN_0;
  wire  _T_7;
  wire [15:0] _GEN_1;
  wire  _T_8;
  assign _T_1 = io_d_in[15:0];
  assign _T_2 = io_d_in[31:16];
  assign _T_3 = io_d_in[47:32];
  assign _T_4 = io_d_in[63:48];
  assign _T_5 = _T_1 > _T_2;
  assign _GEN_0 = _T_5 ? _T_1 : _T_2;
  assign _T_7 = _T_3 > _T_4;
  assign _GEN_1 = _T_7 ? _T_3 : _T_4;
  assign _T_8 = _GEN_0 > _GEN_1;
  assign io_q = _T_8 ? _GEN_0 : _GEN_1;
  assign io_v = io_rdy;
endmodule
module MaxPool1(
  input         clock,
  input         reset,
  input  [15:0] io_d_in,
  input         io_rdy,
  output [15:0] io_d_out,
  output        io_v
);
  wire [63:0] maxpool_io_d_in;
  wire  maxpool_io_rdy;
  wire [15:0] maxpool_io_q;
  wire  maxpool_io_v;
  reg [63:0] pool;
  reg [63:0] _RAND_0;
  reg [2:0] counter;
  reg [31:0] _RAND_1;
  wire  _T;
  wire [3:0] _T_1;
  wire [4:0] _GEN_5;
  wire [7:0] _T_2;
  wire [270:0] _GEN_6;
  wire [270:0] _T_3;
  wire [270:0] _GEN_7;
  wire [271:0] _T_4;
  wire [3:0] _GEN_0;
  wire [3:0] _GEN_2;
  MaxPool maxpool (
    .io_d_in(maxpool_io_d_in),
    .io_rdy(maxpool_io_rdy),
    .io_q(maxpool_io_q),
    .io_v(maxpool_io_v)
  );
  assign _T = counter == 3'h4;
  assign _T_1 = counter + 3'h1;
  assign _GEN_5 = {{2'd0}, counter};
  assign _T_2 = 5'h10 * _GEN_5;
  assign _GEN_6 = {{255'd0}, io_d_in};
  assign _T_3 = _GEN_6 << _T_2;
  assign _GEN_7 = {{207'd0}, pool};
  assign _T_4 = _GEN_7 + _T_3;
  assign _GEN_0 = io_rdy ? _T_1 : {{1'd0}, counter};
  assign _GEN_2 = _T ? 4'h0 : _GEN_0;
  assign io_d_out = maxpool_io_q;
  assign io_v = maxpool_io_v;
  assign maxpool_io_d_in = pool;
  assign maxpool_io_rdy = counter == 3'h4;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pool = _RAND_0[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  counter = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pool <= 64'h0;
    end else if (_T) begin
      pool <= 64'h0;
    end else if (io_rdy) begin
      pool <= _T_4[63:0];
    end
    if (reset) begin
      counter <= 3'h0;
    end else begin
      counter <= _GEN_2[2:0];
    end
  end
endmodule
module Tile(
  input          clock,
  input          reset,
  input  [399:0] io_d_in,
  input  [399:0] io_w_in_0,
  input  [399:0] io_w_in_1,
  input  [399:0] io_w_in_2,
  input  [399:0] io_w_in_3,
  input  [399:0] io_w_in_4,
  input  [399:0] io_w_in_5,
  input  [95:0]  io_bias,
  input          io_rdy,
  output         io_v,
  output [15:0]  io_d_out_0,
  output [15:0]  io_d_out_1,
  output [15:0]  io_d_out_2,
  output [15:0]  io_d_out_3,
  output [15:0]  io_d_out_4,
  output [15:0]  io_d_out_5,
  output         io_pool_v
);
  wire  convc1_clock;
  wire  convc1_reset;
  wire [399:0] convc1_io_d_in;
  wire [399:0] convc1_io_w_in_0;
  wire [399:0] convc1_io_w_in_1;
  wire [399:0] convc1_io_w_in_2;
  wire [399:0] convc1_io_w_in_3;
  wire [399:0] convc1_io_w_in_4;
  wire [399:0] convc1_io_w_in_5;
  wire [95:0] convc1_io_bias;
  wire  convc1_io_rdy;
  wire [15:0] convc1_io_d_out_0;
  wire [15:0] convc1_io_d_out_1;
  wire [15:0] convc1_io_d_out_2;
  wire [15:0] convc1_io_d_out_3;
  wire [15:0] convc1_io_d_out_4;
  wire [15:0] convc1_io_d_out_5;
  wire  convc1_io_v;
  wire  _T_clock;
  wire  _T_reset;
  wire [15:0] _T_io_d_in;
  wire  _T_io_rdy;
  wire [15:0] _T_io_d_out;
  wire  _T_io_v;
  wire  _T_1_clock;
  wire  _T_1_reset;
  wire [15:0] _T_1_io_d_in;
  wire  _T_1_io_rdy;
  wire [15:0] _T_1_io_d_out;
  wire  _T_1_io_v;
  wire  _T_2_clock;
  wire  _T_2_reset;
  wire [15:0] _T_2_io_d_in;
  wire  _T_2_io_rdy;
  wire [15:0] _T_2_io_d_out;
  wire  _T_2_io_v;
  wire  _T_3_clock;
  wire  _T_3_reset;
  wire [15:0] _T_3_io_d_in;
  wire  _T_3_io_rdy;
  wire [15:0] _T_3_io_d_out;
  wire  _T_3_io_v;
  wire  _T_4_clock;
  wire  _T_4_reset;
  wire [15:0] _T_4_io_d_in;
  wire  _T_4_io_rdy;
  wire [15:0] _T_4_io_d_out;
  wire  _T_4_io_v;
  wire  _T_5_clock;
  wire  _T_5_reset;
  wire [15:0] _T_5_io_d_in;
  wire  _T_5_io_rdy;
  wire [15:0] _T_5_io_d_out;
  wire  _T_5_io_v;
  wire  _T_6;
  wire  _T_7;
  wire  _T_8;
  wire  _T_9;
  ConvC1 convc1 (
    .clock(convc1_clock),
    .reset(convc1_reset),
    .io_d_in(convc1_io_d_in),
    .io_w_in_0(convc1_io_w_in_0),
    .io_w_in_1(convc1_io_w_in_1),
    .io_w_in_2(convc1_io_w_in_2),
    .io_w_in_3(convc1_io_w_in_3),
    .io_w_in_4(convc1_io_w_in_4),
    .io_w_in_5(convc1_io_w_in_5),
    .io_bias(convc1_io_bias),
    .io_rdy(convc1_io_rdy),
    .io_d_out_0(convc1_io_d_out_0),
    .io_d_out_1(convc1_io_d_out_1),
    .io_d_out_2(convc1_io_d_out_2),
    .io_d_out_3(convc1_io_d_out_3),
    .io_d_out_4(convc1_io_d_out_4),
    .io_d_out_5(convc1_io_d_out_5),
    .io_v(convc1_io_v)
  );
  MaxPool1 _T (
    .clock(_T_clock),
    .reset(_T_reset),
    .io_d_in(_T_io_d_in),
    .io_rdy(_T_io_rdy),
    .io_d_out(_T_io_d_out),
    .io_v(_T_io_v)
  );
  MaxPool1 _T_1 (
    .clock(_T_1_clock),
    .reset(_T_1_reset),
    .io_d_in(_T_1_io_d_in),
    .io_rdy(_T_1_io_rdy),
    .io_d_out(_T_1_io_d_out),
    .io_v(_T_1_io_v)
  );
  MaxPool1 _T_2 (
    .clock(_T_2_clock),
    .reset(_T_2_reset),
    .io_d_in(_T_2_io_d_in),
    .io_rdy(_T_2_io_rdy),
    .io_d_out(_T_2_io_d_out),
    .io_v(_T_2_io_v)
  );
  MaxPool1 _T_3 (
    .clock(_T_3_clock),
    .reset(_T_3_reset),
    .io_d_in(_T_3_io_d_in),
    .io_rdy(_T_3_io_rdy),
    .io_d_out(_T_3_io_d_out),
    .io_v(_T_3_io_v)
  );
  MaxPool1 _T_4 (
    .clock(_T_4_clock),
    .reset(_T_4_reset),
    .io_d_in(_T_4_io_d_in),
    .io_rdy(_T_4_io_rdy),
    .io_d_out(_T_4_io_d_out),
    .io_v(_T_4_io_v)
  );
  MaxPool1 _T_5 (
    .clock(_T_5_clock),
    .reset(_T_5_reset),
    .io_d_in(_T_5_io_d_in),
    .io_rdy(_T_5_io_rdy),
    .io_d_out(_T_5_io_d_out),
    .io_v(_T_5_io_v)
  );
  assign _T_6 = _T_io_v & _T_1_io_v;
  assign _T_7 = _T_6 & _T_2_io_v;
  assign _T_8 = _T_7 & _T_3_io_v;
  assign _T_9 = _T_8 & _T_4_io_v;
  assign io_v = convc1_io_v;
  assign io_d_out_0 = _T_io_d_out;
  assign io_d_out_1 = _T_1_io_d_out;
  assign io_d_out_2 = _T_2_io_d_out;
  assign io_d_out_3 = _T_3_io_d_out;
  assign io_d_out_4 = _T_4_io_d_out;
  assign io_d_out_5 = _T_5_io_d_out;
  assign io_pool_v = _T_9 & _T_5_io_v;
  assign convc1_clock = clock;
  assign convc1_reset = reset;
  assign convc1_io_d_in = io_d_in;
  assign convc1_io_w_in_0 = io_w_in_0;
  assign convc1_io_w_in_1 = io_w_in_1;
  assign convc1_io_w_in_2 = io_w_in_2;
  assign convc1_io_w_in_3 = io_w_in_3;
  assign convc1_io_w_in_4 = io_w_in_4;
  assign convc1_io_w_in_5 = io_w_in_5;
  assign convc1_io_bias = io_bias;
  assign convc1_io_rdy = io_rdy;
  assign _T_clock = clock;
  assign _T_reset = reset;
  assign _T_io_d_in = convc1_io_d_out_0;
  assign _T_io_rdy = convc1_io_v;
  assign _T_1_clock = clock;
  assign _T_1_reset = reset;
  assign _T_1_io_d_in = convc1_io_d_out_1;
  assign _T_1_io_rdy = convc1_io_v;
  assign _T_2_clock = clock;
  assign _T_2_reset = reset;
  assign _T_2_io_d_in = convc1_io_d_out_2;
  assign _T_2_io_rdy = convc1_io_v;
  assign _T_3_clock = clock;
  assign _T_3_reset = reset;
  assign _T_3_io_d_in = convc1_io_d_out_3;
  assign _T_3_io_rdy = convc1_io_v;
  assign _T_4_clock = clock;
  assign _T_4_reset = reset;
  assign _T_4_io_d_in = convc1_io_d_out_4;
  assign _T_4_io_rdy = convc1_io_v;
  assign _T_5_clock = clock;
  assign _T_5_reset = reset;
  assign _T_5_io_d_in = convc1_io_d_out_5;
  assign _T_5_io_rdy = convc1_io_v;
endmodule
module ShiftRegister(
  input          clock,
  input          reset,
  input  [15:0]  io_d_in,
  input          io_en,
  output [399:0] io_d_out
);
  reg [15:0] _T;
  reg [31:0] _RAND_0;
  reg [15:0] _T_1;
  reg [31:0] _RAND_1;
  reg [15:0] _T_2;
  reg [31:0] _RAND_2;
  reg [15:0] _T_3;
  reg [31:0] _RAND_3;
  reg [15:0] _T_4;
  reg [31:0] _RAND_4;
  reg [15:0] _T_5;
  reg [31:0] _RAND_5;
  reg [15:0] _T_6;
  reg [31:0] _RAND_6;
  reg [15:0] _T_7;
  reg [31:0] _RAND_7;
  reg [15:0] _T_8;
  reg [31:0] _RAND_8;
  reg [15:0] _T_9;
  reg [31:0] _RAND_9;
  reg [15:0] _T_10;
  reg [31:0] _RAND_10;
  reg [15:0] _T_11;
  reg [31:0] _RAND_11;
  reg [15:0] _T_12;
  reg [31:0] _RAND_12;
  reg [15:0] _T_13;
  reg [31:0] _RAND_13;
  reg [15:0] _T_14;
  reg [31:0] _RAND_14;
  reg [15:0] _T_15;
  reg [31:0] _RAND_15;
  reg [15:0] _T_16;
  reg [31:0] _RAND_16;
  reg [15:0] _T_17;
  reg [31:0] _RAND_17;
  reg [15:0] _T_18;
  reg [31:0] _RAND_18;
  reg [15:0] _T_19;
  reg [31:0] _RAND_19;
  reg [15:0] _T_20;
  reg [31:0] _RAND_20;
  reg [15:0] _T_21;
  reg [31:0] _RAND_21;
  reg [15:0] _T_22;
  reg [31:0] _RAND_22;
  reg [15:0] _T_23;
  reg [31:0] _RAND_23;
  reg [15:0] _T_24;
  reg [31:0] _RAND_24;
  wire [95:0] _T_34;
  wire [191:0] _T_35;
  wire [111:0] _T_46;
  wire [207:0] _T_47;
  assign _T_34 = {_T_6,_T_7,_T_8,_T_9,_T_10,_T_11};
  assign _T_35 = {_T,_T_1,_T_2,_T_3,_T_4,_T_5,_T_34};
  assign _T_46 = {_T_18,_T_19,_T_20,_T_21,_T_22,_T_23,_T_24};
  assign _T_47 = {_T_12,_T_13,_T_14,_T_15,_T_16,_T_17,_T_46};
  assign io_d_out = {_T_35,_T_47};
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_6 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_7 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_8 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_9 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_10 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_11 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_12 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_13 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_14 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_15 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_16 = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_17 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_18 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_19 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_20 = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_21 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_22 = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_23 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_24 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T <= 16'h0;
    end else if (io_en) begin
      _T <= io_d_in;
    end
    if (reset) begin
      _T_1 <= 16'h0;
    end else if (io_en) begin
      _T_1 <= _T;
    end
    if (reset) begin
      _T_2 <= 16'h0;
    end else if (io_en) begin
      _T_2 <= _T_1;
    end
    if (reset) begin
      _T_3 <= 16'h0;
    end else if (io_en) begin
      _T_3 <= _T_2;
    end
    if (reset) begin
      _T_4 <= 16'h0;
    end else if (io_en) begin
      _T_4 <= _T_3;
    end
    if (reset) begin
      _T_5 <= 16'h0;
    end else if (io_en) begin
      _T_5 <= _T_4;
    end
    if (reset) begin
      _T_6 <= 16'h0;
    end else if (io_en) begin
      _T_6 <= _T_5;
    end
    if (reset) begin
      _T_7 <= 16'h0;
    end else if (io_en) begin
      _T_7 <= _T_6;
    end
    if (reset) begin
      _T_8 <= 16'h0;
    end else if (io_en) begin
      _T_8 <= _T_7;
    end
    if (reset) begin
      _T_9 <= 16'h0;
    end else if (io_en) begin
      _T_9 <= _T_8;
    end
    if (reset) begin
      _T_10 <= 16'h0;
    end else if (io_en) begin
      _T_10 <= _T_9;
    end
    if (reset) begin
      _T_11 <= 16'h0;
    end else if (io_en) begin
      _T_11 <= _T_10;
    end
    if (reset) begin
      _T_12 <= 16'h0;
    end else if (io_en) begin
      _T_12 <= _T_11;
    end
    if (reset) begin
      _T_13 <= 16'h0;
    end else if (io_en) begin
      _T_13 <= _T_12;
    end
    if (reset) begin
      _T_14 <= 16'h0;
    end else if (io_en) begin
      _T_14 <= _T_13;
    end
    if (reset) begin
      _T_15 <= 16'h0;
    end else if (io_en) begin
      _T_15 <= _T_14;
    end
    if (reset) begin
      _T_16 <= 16'h0;
    end else if (io_en) begin
      _T_16 <= _T_15;
    end
    if (reset) begin
      _T_17 <= 16'h0;
    end else if (io_en) begin
      _T_17 <= _T_16;
    end
    if (reset) begin
      _T_18 <= 16'h0;
    end else if (io_en) begin
      _T_18 <= _T_17;
    end
    if (reset) begin
      _T_19 <= 16'h0;
    end else if (io_en) begin
      _T_19 <= _T_18;
    end
    if (reset) begin
      _T_20 <= 16'h0;
    end else if (io_en) begin
      _T_20 <= _T_19;
    end
    if (reset) begin
      _T_21 <= 16'h0;
    end else if (io_en) begin
      _T_21 <= _T_20;
    end
    if (reset) begin
      _T_22 <= 16'h0;
    end else if (io_en) begin
      _T_22 <= _T_21;
    end
    if (reset) begin
      _T_23 <= 16'h0;
    end else if (io_en) begin
      _T_23 <= _T_22;
    end
    if (reset) begin
      _T_24 <= 16'h0;
    end else if (io_en) begin
      _T_24 <= _T_23;
    end
  end
endmodule
module ConvC3(
  input          clock,
  input          reset,
  input  [399:0] io_d_in,
  input  [399:0] io_w_in_0,
  input  [399:0] io_w_in_1,
  input  [399:0] io_w_in_2,
  input  [399:0] io_w_in_3,
  input  [399:0] io_w_in_4,
  input  [399:0] io_w_in_5,
  input  [399:0] io_w_in_6,
  input  [399:0] io_w_in_7,
  input  [399:0] io_w_in_8,
  input  [399:0] io_w_in_9,
  input  [399:0] io_w_in_10,
  input  [399:0] io_w_in_11,
  input  [399:0] io_w_in_12,
  input  [399:0] io_w_in_13,
  input  [399:0] io_w_in_14,
  input  [399:0] io_w_in_15,
  input          io_rdy,
  output [15:0]  io_d_out_0,
  output [15:0]  io_d_out_1,
  output [15:0]  io_d_out_2,
  output [15:0]  io_d_out_3,
  output [15:0]  io_d_out_4,
  output [15:0]  io_d_out_5,
  output [15:0]  io_d_out_6,
  output [15:0]  io_d_out_7,
  output [15:0]  io_d_out_8,
  output [15:0]  io_d_out_9,
  output [15:0]  io_d_out_10,
  output [15:0]  io_d_out_11,
  output [15:0]  io_d_out_12,
  output [15:0]  io_d_out_13,
  output [15:0]  io_d_out_14,
  output [15:0]  io_d_out_15,
  output         io_v
);
  wire  _T_clock;
  wire  _T_reset;
  wire [399:0] _T_io_d_in;
  wire [399:0] _T_io_w;
  wire  _T_io_rdy;
  wire [15:0] _T_io_bias;
  wire [15:0] _T_io_d_out;
  wire  _T_io_v;
  wire  _T_1_clock;
  wire  _T_1_reset;
  wire [399:0] _T_1_io_d_in;
  wire [399:0] _T_1_io_w;
  wire  _T_1_io_rdy;
  wire [15:0] _T_1_io_bias;
  wire [15:0] _T_1_io_d_out;
  wire  _T_1_io_v;
  wire  _T_2_clock;
  wire  _T_2_reset;
  wire [399:0] _T_2_io_d_in;
  wire [399:0] _T_2_io_w;
  wire  _T_2_io_rdy;
  wire [15:0] _T_2_io_bias;
  wire [15:0] _T_2_io_d_out;
  wire  _T_2_io_v;
  wire  _T_3_clock;
  wire  _T_3_reset;
  wire [399:0] _T_3_io_d_in;
  wire [399:0] _T_3_io_w;
  wire  _T_3_io_rdy;
  wire [15:0] _T_3_io_bias;
  wire [15:0] _T_3_io_d_out;
  wire  _T_3_io_v;
  wire  _T_4_clock;
  wire  _T_4_reset;
  wire [399:0] _T_4_io_d_in;
  wire [399:0] _T_4_io_w;
  wire  _T_4_io_rdy;
  wire [15:0] _T_4_io_bias;
  wire [15:0] _T_4_io_d_out;
  wire  _T_4_io_v;
  wire  _T_5_clock;
  wire  _T_5_reset;
  wire [399:0] _T_5_io_d_in;
  wire [399:0] _T_5_io_w;
  wire  _T_5_io_rdy;
  wire [15:0] _T_5_io_bias;
  wire [15:0] _T_5_io_d_out;
  wire  _T_5_io_v;
  wire  _T_6_clock;
  wire  _T_6_reset;
  wire [399:0] _T_6_io_d_in;
  wire [399:0] _T_6_io_w;
  wire  _T_6_io_rdy;
  wire [15:0] _T_6_io_bias;
  wire [15:0] _T_6_io_d_out;
  wire  _T_6_io_v;
  wire  _T_7_clock;
  wire  _T_7_reset;
  wire [399:0] _T_7_io_d_in;
  wire [399:0] _T_7_io_w;
  wire  _T_7_io_rdy;
  wire [15:0] _T_7_io_bias;
  wire [15:0] _T_7_io_d_out;
  wire  _T_7_io_v;
  wire  _T_8_clock;
  wire  _T_8_reset;
  wire [399:0] _T_8_io_d_in;
  wire [399:0] _T_8_io_w;
  wire  _T_8_io_rdy;
  wire [15:0] _T_8_io_bias;
  wire [15:0] _T_8_io_d_out;
  wire  _T_8_io_v;
  wire  _T_9_clock;
  wire  _T_9_reset;
  wire [399:0] _T_9_io_d_in;
  wire [399:0] _T_9_io_w;
  wire  _T_9_io_rdy;
  wire [15:0] _T_9_io_bias;
  wire [15:0] _T_9_io_d_out;
  wire  _T_9_io_v;
  wire  _T_10_clock;
  wire  _T_10_reset;
  wire [399:0] _T_10_io_d_in;
  wire [399:0] _T_10_io_w;
  wire  _T_10_io_rdy;
  wire [15:0] _T_10_io_bias;
  wire [15:0] _T_10_io_d_out;
  wire  _T_10_io_v;
  wire  _T_11_clock;
  wire  _T_11_reset;
  wire [399:0] _T_11_io_d_in;
  wire [399:0] _T_11_io_w;
  wire  _T_11_io_rdy;
  wire [15:0] _T_11_io_bias;
  wire [15:0] _T_11_io_d_out;
  wire  _T_11_io_v;
  wire  _T_12_clock;
  wire  _T_12_reset;
  wire [399:0] _T_12_io_d_in;
  wire [399:0] _T_12_io_w;
  wire  _T_12_io_rdy;
  wire [15:0] _T_12_io_bias;
  wire [15:0] _T_12_io_d_out;
  wire  _T_12_io_v;
  wire  _T_13_clock;
  wire  _T_13_reset;
  wire [399:0] _T_13_io_d_in;
  wire [399:0] _T_13_io_w;
  wire  _T_13_io_rdy;
  wire [15:0] _T_13_io_bias;
  wire [15:0] _T_13_io_d_out;
  wire  _T_13_io_v;
  wire  _T_14_clock;
  wire  _T_14_reset;
  wire [399:0] _T_14_io_d_in;
  wire [399:0] _T_14_io_w;
  wire  _T_14_io_rdy;
  wire [15:0] _T_14_io_bias;
  wire [15:0] _T_14_io_d_out;
  wire  _T_14_io_v;
  wire  _T_15_clock;
  wire  _T_15_reset;
  wire [399:0] _T_15_io_d_in;
  wire [399:0] _T_15_io_w;
  wire  _T_15_io_rdy;
  wire [15:0] _T_15_io_bias;
  wire [15:0] _T_15_io_d_out;
  wire  _T_15_io_v;
  wire  _T_16;
  wire  _T_17;
  wire  _T_18;
  wire  _T_19;
  wire  _T_20;
  wire  _T_21;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_26;
  wire  _T_27;
  wire  _T_28;
  wire  _T_29;
  Node _T (
    .clock(_T_clock),
    .reset(_T_reset),
    .io_d_in(_T_io_d_in),
    .io_w(_T_io_w),
    .io_rdy(_T_io_rdy),
    .io_bias(_T_io_bias),
    .io_d_out(_T_io_d_out),
    .io_v(_T_io_v)
  );
  Node _T_1 (
    .clock(_T_1_clock),
    .reset(_T_1_reset),
    .io_d_in(_T_1_io_d_in),
    .io_w(_T_1_io_w),
    .io_rdy(_T_1_io_rdy),
    .io_bias(_T_1_io_bias),
    .io_d_out(_T_1_io_d_out),
    .io_v(_T_1_io_v)
  );
  Node _T_2 (
    .clock(_T_2_clock),
    .reset(_T_2_reset),
    .io_d_in(_T_2_io_d_in),
    .io_w(_T_2_io_w),
    .io_rdy(_T_2_io_rdy),
    .io_bias(_T_2_io_bias),
    .io_d_out(_T_2_io_d_out),
    .io_v(_T_2_io_v)
  );
  Node _T_3 (
    .clock(_T_3_clock),
    .reset(_T_3_reset),
    .io_d_in(_T_3_io_d_in),
    .io_w(_T_3_io_w),
    .io_rdy(_T_3_io_rdy),
    .io_bias(_T_3_io_bias),
    .io_d_out(_T_3_io_d_out),
    .io_v(_T_3_io_v)
  );
  Node _T_4 (
    .clock(_T_4_clock),
    .reset(_T_4_reset),
    .io_d_in(_T_4_io_d_in),
    .io_w(_T_4_io_w),
    .io_rdy(_T_4_io_rdy),
    .io_bias(_T_4_io_bias),
    .io_d_out(_T_4_io_d_out),
    .io_v(_T_4_io_v)
  );
  Node _T_5 (
    .clock(_T_5_clock),
    .reset(_T_5_reset),
    .io_d_in(_T_5_io_d_in),
    .io_w(_T_5_io_w),
    .io_rdy(_T_5_io_rdy),
    .io_bias(_T_5_io_bias),
    .io_d_out(_T_5_io_d_out),
    .io_v(_T_5_io_v)
  );
  Node _T_6 (
    .clock(_T_6_clock),
    .reset(_T_6_reset),
    .io_d_in(_T_6_io_d_in),
    .io_w(_T_6_io_w),
    .io_rdy(_T_6_io_rdy),
    .io_bias(_T_6_io_bias),
    .io_d_out(_T_6_io_d_out),
    .io_v(_T_6_io_v)
  );
  Node _T_7 (
    .clock(_T_7_clock),
    .reset(_T_7_reset),
    .io_d_in(_T_7_io_d_in),
    .io_w(_T_7_io_w),
    .io_rdy(_T_7_io_rdy),
    .io_bias(_T_7_io_bias),
    .io_d_out(_T_7_io_d_out),
    .io_v(_T_7_io_v)
  );
  Node _T_8 (
    .clock(_T_8_clock),
    .reset(_T_8_reset),
    .io_d_in(_T_8_io_d_in),
    .io_w(_T_8_io_w),
    .io_rdy(_T_8_io_rdy),
    .io_bias(_T_8_io_bias),
    .io_d_out(_T_8_io_d_out),
    .io_v(_T_8_io_v)
  );
  Node _T_9 (
    .clock(_T_9_clock),
    .reset(_T_9_reset),
    .io_d_in(_T_9_io_d_in),
    .io_w(_T_9_io_w),
    .io_rdy(_T_9_io_rdy),
    .io_bias(_T_9_io_bias),
    .io_d_out(_T_9_io_d_out),
    .io_v(_T_9_io_v)
  );
  Node _T_10 (
    .clock(_T_10_clock),
    .reset(_T_10_reset),
    .io_d_in(_T_10_io_d_in),
    .io_w(_T_10_io_w),
    .io_rdy(_T_10_io_rdy),
    .io_bias(_T_10_io_bias),
    .io_d_out(_T_10_io_d_out),
    .io_v(_T_10_io_v)
  );
  Node _T_11 (
    .clock(_T_11_clock),
    .reset(_T_11_reset),
    .io_d_in(_T_11_io_d_in),
    .io_w(_T_11_io_w),
    .io_rdy(_T_11_io_rdy),
    .io_bias(_T_11_io_bias),
    .io_d_out(_T_11_io_d_out),
    .io_v(_T_11_io_v)
  );
  Node _T_12 (
    .clock(_T_12_clock),
    .reset(_T_12_reset),
    .io_d_in(_T_12_io_d_in),
    .io_w(_T_12_io_w),
    .io_rdy(_T_12_io_rdy),
    .io_bias(_T_12_io_bias),
    .io_d_out(_T_12_io_d_out),
    .io_v(_T_12_io_v)
  );
  Node _T_13 (
    .clock(_T_13_clock),
    .reset(_T_13_reset),
    .io_d_in(_T_13_io_d_in),
    .io_w(_T_13_io_w),
    .io_rdy(_T_13_io_rdy),
    .io_bias(_T_13_io_bias),
    .io_d_out(_T_13_io_d_out),
    .io_v(_T_13_io_v)
  );
  Node _T_14 (
    .clock(_T_14_clock),
    .reset(_T_14_reset),
    .io_d_in(_T_14_io_d_in),
    .io_w(_T_14_io_w),
    .io_rdy(_T_14_io_rdy),
    .io_bias(_T_14_io_bias),
    .io_d_out(_T_14_io_d_out),
    .io_v(_T_14_io_v)
  );
  Node _T_15 (
    .clock(_T_15_clock),
    .reset(_T_15_reset),
    .io_d_in(_T_15_io_d_in),
    .io_w(_T_15_io_w),
    .io_rdy(_T_15_io_rdy),
    .io_bias(_T_15_io_bias),
    .io_d_out(_T_15_io_d_out),
    .io_v(_T_15_io_v)
  );
  assign _T_16 = _T_io_v & _T_1_io_v;
  assign _T_17 = _T_16 & _T_2_io_v;
  assign _T_18 = _T_17 & _T_3_io_v;
  assign _T_19 = _T_18 & _T_4_io_v;
  assign _T_20 = _T_19 & _T_5_io_v;
  assign _T_21 = _T_20 & _T_6_io_v;
  assign _T_22 = _T_21 & _T_7_io_v;
  assign _T_23 = _T_22 & _T_8_io_v;
  assign _T_24 = _T_23 & _T_9_io_v;
  assign _T_25 = _T_24 & _T_10_io_v;
  assign _T_26 = _T_25 & _T_11_io_v;
  assign _T_27 = _T_26 & _T_12_io_v;
  assign _T_28 = _T_27 & _T_13_io_v;
  assign _T_29 = _T_28 & _T_14_io_v;
  assign io_d_out_0 = _T_io_d_out;
  assign io_d_out_1 = _T_1_io_d_out;
  assign io_d_out_2 = _T_2_io_d_out;
  assign io_d_out_3 = _T_3_io_d_out;
  assign io_d_out_4 = _T_4_io_d_out;
  assign io_d_out_5 = _T_5_io_d_out;
  assign io_d_out_6 = _T_6_io_d_out;
  assign io_d_out_7 = _T_7_io_d_out;
  assign io_d_out_8 = _T_8_io_d_out;
  assign io_d_out_9 = _T_9_io_d_out;
  assign io_d_out_10 = _T_10_io_d_out;
  assign io_d_out_11 = _T_11_io_d_out;
  assign io_d_out_12 = _T_12_io_d_out;
  assign io_d_out_13 = _T_13_io_d_out;
  assign io_d_out_14 = _T_14_io_d_out;
  assign io_d_out_15 = _T_15_io_d_out;
  assign io_v = _T_29 & _T_15_io_v;
  assign _T_clock = clock;
  assign _T_reset = reset;
  assign _T_io_d_in = io_d_in;
  assign _T_io_w = io_w_in_0;
  assign _T_io_rdy = io_rdy;
  assign _T_io_bias = 16'h0;
  assign _T_1_clock = clock;
  assign _T_1_reset = reset;
  assign _T_1_io_d_in = io_d_in;
  assign _T_1_io_w = io_w_in_1;
  assign _T_1_io_rdy = io_rdy;
  assign _T_1_io_bias = 16'h0;
  assign _T_2_clock = clock;
  assign _T_2_reset = reset;
  assign _T_2_io_d_in = io_d_in;
  assign _T_2_io_w = io_w_in_2;
  assign _T_2_io_rdy = io_rdy;
  assign _T_2_io_bias = 16'h0;
  assign _T_3_clock = clock;
  assign _T_3_reset = reset;
  assign _T_3_io_d_in = io_d_in;
  assign _T_3_io_w = io_w_in_3;
  assign _T_3_io_rdy = io_rdy;
  assign _T_3_io_bias = 16'h0;
  assign _T_4_clock = clock;
  assign _T_4_reset = reset;
  assign _T_4_io_d_in = io_d_in;
  assign _T_4_io_w = io_w_in_4;
  assign _T_4_io_rdy = io_rdy;
  assign _T_4_io_bias = 16'h0;
  assign _T_5_clock = clock;
  assign _T_5_reset = reset;
  assign _T_5_io_d_in = io_d_in;
  assign _T_5_io_w = io_w_in_5;
  assign _T_5_io_rdy = io_rdy;
  assign _T_5_io_bias = 16'h0;
  assign _T_6_clock = clock;
  assign _T_6_reset = reset;
  assign _T_6_io_d_in = io_d_in;
  assign _T_6_io_w = io_w_in_6;
  assign _T_6_io_rdy = io_rdy;
  assign _T_6_io_bias = 16'h0;
  assign _T_7_clock = clock;
  assign _T_7_reset = reset;
  assign _T_7_io_d_in = io_d_in;
  assign _T_7_io_w = io_w_in_7;
  assign _T_7_io_rdy = io_rdy;
  assign _T_7_io_bias = 16'h0;
  assign _T_8_clock = clock;
  assign _T_8_reset = reset;
  assign _T_8_io_d_in = io_d_in;
  assign _T_8_io_w = io_w_in_8;
  assign _T_8_io_rdy = io_rdy;
  assign _T_8_io_bias = 16'h0;
  assign _T_9_clock = clock;
  assign _T_9_reset = reset;
  assign _T_9_io_d_in = io_d_in;
  assign _T_9_io_w = io_w_in_9;
  assign _T_9_io_rdy = io_rdy;
  assign _T_9_io_bias = 16'h0;
  assign _T_10_clock = clock;
  assign _T_10_reset = reset;
  assign _T_10_io_d_in = io_d_in;
  assign _T_10_io_w = io_w_in_10;
  assign _T_10_io_rdy = io_rdy;
  assign _T_10_io_bias = 16'h0;
  assign _T_11_clock = clock;
  assign _T_11_reset = reset;
  assign _T_11_io_d_in = io_d_in;
  assign _T_11_io_w = io_w_in_11;
  assign _T_11_io_rdy = io_rdy;
  assign _T_11_io_bias = 16'h0;
  assign _T_12_clock = clock;
  assign _T_12_reset = reset;
  assign _T_12_io_d_in = io_d_in;
  assign _T_12_io_w = io_w_in_12;
  assign _T_12_io_rdy = io_rdy;
  assign _T_12_io_bias = 16'h0;
  assign _T_13_clock = clock;
  assign _T_13_reset = reset;
  assign _T_13_io_d_in = io_d_in;
  assign _T_13_io_w = io_w_in_13;
  assign _T_13_io_rdy = io_rdy;
  assign _T_13_io_bias = 16'h0;
  assign _T_14_clock = clock;
  assign _T_14_reset = reset;
  assign _T_14_io_d_in = io_d_in;
  assign _T_14_io_w = io_w_in_14;
  assign _T_14_io_rdy = io_rdy;
  assign _T_14_io_bias = 16'h0;
  assign _T_15_clock = clock;
  assign _T_15_reset = reset;
  assign _T_15_io_d_in = io_d_in;
  assign _T_15_io_w = io_w_in_15;
  assign _T_15_io_rdy = io_rdy;
  assign _T_15_io_bias = 16'h0;
endmodule
module Tile2(
  input         clock,
  input         reset,
  input  [15:0] io_d_in_0,
  input  [15:0] io_d_in_1,
  input  [15:0] io_d_in_2,
  input  [15:0] io_d_in_3,
  input  [15:0] io_d_in_4,
  input  [15:0] io_d_in_5,
  input         io_rdy,
  output        io_c3_v,
  output [15:0] io_d_out_0,
  output [15:0] io_d_out_1,
  output [15:0] io_d_out_2,
  output [15:0] io_d_out_3,
  output [15:0] io_d_out_4,
  output [15:0] io_d_out_5,
  output [15:0] io_d_out_6,
  output [15:0] io_d_out_7,
  output [15:0] io_d_out_8,
  output [15:0] io_d_out_9,
  output [15:0] io_d_out_10,
  output [15:0] io_d_out_11,
  output [15:0] io_d_out_12,
  output [15:0] io_d_out_13,
  output [15:0] io_d_out_14,
  output [15:0] io_d_out_15
);
  wire  _T_clock;
  wire  _T_reset;
  wire [15:0] _T_io_d_in;
  wire  _T_io_en;
  wire [399:0] _T_io_d_out;
  wire  _T_1_clock;
  wire  _T_1_reset;
  wire [399:0] _T_1_io_d_in;
  wire [399:0] _T_1_io_w_in_0;
  wire [399:0] _T_1_io_w_in_1;
  wire [399:0] _T_1_io_w_in_2;
  wire [399:0] _T_1_io_w_in_3;
  wire [399:0] _T_1_io_w_in_4;
  wire [399:0] _T_1_io_w_in_5;
  wire [399:0] _T_1_io_w_in_6;
  wire [399:0] _T_1_io_w_in_7;
  wire [399:0] _T_1_io_w_in_8;
  wire [399:0] _T_1_io_w_in_9;
  wire [399:0] _T_1_io_w_in_10;
  wire [399:0] _T_1_io_w_in_11;
  wire [399:0] _T_1_io_w_in_12;
  wire [399:0] _T_1_io_w_in_13;
  wire [399:0] _T_1_io_w_in_14;
  wire [399:0] _T_1_io_w_in_15;
  wire  _T_1_io_rdy;
  wire [15:0] _T_1_io_d_out_0;
  wire [15:0] _T_1_io_d_out_1;
  wire [15:0] _T_1_io_d_out_2;
  wire [15:0] _T_1_io_d_out_3;
  wire [15:0] _T_1_io_d_out_4;
  wire [15:0] _T_1_io_d_out_5;
  wire [15:0] _T_1_io_d_out_6;
  wire [15:0] _T_1_io_d_out_7;
  wire [15:0] _T_1_io_d_out_8;
  wire [15:0] _T_1_io_d_out_9;
  wire [15:0] _T_1_io_d_out_10;
  wire [15:0] _T_1_io_d_out_11;
  wire [15:0] _T_1_io_d_out_12;
  wire [15:0] _T_1_io_d_out_13;
  wire [15:0] _T_1_io_d_out_14;
  wire [15:0] _T_1_io_d_out_15;
  wire  _T_1_io_v;
  wire  _T_2_clock;
  wire  _T_2_reset;
  wire [15:0] _T_2_io_d_in;
  wire  _T_2_io_en;
  wire [399:0] _T_2_io_d_out;
  wire  _T_3_clock;
  wire  _T_3_reset;
  wire [399:0] _T_3_io_d_in;
  wire [399:0] _T_3_io_w_in_0;
  wire [399:0] _T_3_io_w_in_1;
  wire [399:0] _T_3_io_w_in_2;
  wire [399:0] _T_3_io_w_in_3;
  wire [399:0] _T_3_io_w_in_4;
  wire [399:0] _T_3_io_w_in_5;
  wire [399:0] _T_3_io_w_in_6;
  wire [399:0] _T_3_io_w_in_7;
  wire [399:0] _T_3_io_w_in_8;
  wire [399:0] _T_3_io_w_in_9;
  wire [399:0] _T_3_io_w_in_10;
  wire [399:0] _T_3_io_w_in_11;
  wire [399:0] _T_3_io_w_in_12;
  wire [399:0] _T_3_io_w_in_13;
  wire [399:0] _T_3_io_w_in_14;
  wire [399:0] _T_3_io_w_in_15;
  wire  _T_3_io_rdy;
  wire [15:0] _T_3_io_d_out_0;
  wire [15:0] _T_3_io_d_out_1;
  wire [15:0] _T_3_io_d_out_2;
  wire [15:0] _T_3_io_d_out_3;
  wire [15:0] _T_3_io_d_out_4;
  wire [15:0] _T_3_io_d_out_5;
  wire [15:0] _T_3_io_d_out_6;
  wire [15:0] _T_3_io_d_out_7;
  wire [15:0] _T_3_io_d_out_8;
  wire [15:0] _T_3_io_d_out_9;
  wire [15:0] _T_3_io_d_out_10;
  wire [15:0] _T_3_io_d_out_11;
  wire [15:0] _T_3_io_d_out_12;
  wire [15:0] _T_3_io_d_out_13;
  wire [15:0] _T_3_io_d_out_14;
  wire [15:0] _T_3_io_d_out_15;
  wire  _T_3_io_v;
  wire  _T_4_clock;
  wire  _T_4_reset;
  wire [15:0] _T_4_io_d_in;
  wire  _T_4_io_en;
  wire [399:0] _T_4_io_d_out;
  wire  _T_5_clock;
  wire  _T_5_reset;
  wire [399:0] _T_5_io_d_in;
  wire [399:0] _T_5_io_w_in_0;
  wire [399:0] _T_5_io_w_in_1;
  wire [399:0] _T_5_io_w_in_2;
  wire [399:0] _T_5_io_w_in_3;
  wire [399:0] _T_5_io_w_in_4;
  wire [399:0] _T_5_io_w_in_5;
  wire [399:0] _T_5_io_w_in_6;
  wire [399:0] _T_5_io_w_in_7;
  wire [399:0] _T_5_io_w_in_8;
  wire [399:0] _T_5_io_w_in_9;
  wire [399:0] _T_5_io_w_in_10;
  wire [399:0] _T_5_io_w_in_11;
  wire [399:0] _T_5_io_w_in_12;
  wire [399:0] _T_5_io_w_in_13;
  wire [399:0] _T_5_io_w_in_14;
  wire [399:0] _T_5_io_w_in_15;
  wire  _T_5_io_rdy;
  wire [15:0] _T_5_io_d_out_0;
  wire [15:0] _T_5_io_d_out_1;
  wire [15:0] _T_5_io_d_out_2;
  wire [15:0] _T_5_io_d_out_3;
  wire [15:0] _T_5_io_d_out_4;
  wire [15:0] _T_5_io_d_out_5;
  wire [15:0] _T_5_io_d_out_6;
  wire [15:0] _T_5_io_d_out_7;
  wire [15:0] _T_5_io_d_out_8;
  wire [15:0] _T_5_io_d_out_9;
  wire [15:0] _T_5_io_d_out_10;
  wire [15:0] _T_5_io_d_out_11;
  wire [15:0] _T_5_io_d_out_12;
  wire [15:0] _T_5_io_d_out_13;
  wire [15:0] _T_5_io_d_out_14;
  wire [15:0] _T_5_io_d_out_15;
  wire  _T_5_io_v;
  wire  _T_6_clock;
  wire  _T_6_reset;
  wire [15:0] _T_6_io_d_in;
  wire  _T_6_io_en;
  wire [399:0] _T_6_io_d_out;
  wire  _T_7_clock;
  wire  _T_7_reset;
  wire [399:0] _T_7_io_d_in;
  wire [399:0] _T_7_io_w_in_0;
  wire [399:0] _T_7_io_w_in_1;
  wire [399:0] _T_7_io_w_in_2;
  wire [399:0] _T_7_io_w_in_3;
  wire [399:0] _T_7_io_w_in_4;
  wire [399:0] _T_7_io_w_in_5;
  wire [399:0] _T_7_io_w_in_6;
  wire [399:0] _T_7_io_w_in_7;
  wire [399:0] _T_7_io_w_in_8;
  wire [399:0] _T_7_io_w_in_9;
  wire [399:0] _T_7_io_w_in_10;
  wire [399:0] _T_7_io_w_in_11;
  wire [399:0] _T_7_io_w_in_12;
  wire [399:0] _T_7_io_w_in_13;
  wire [399:0] _T_7_io_w_in_14;
  wire [399:0] _T_7_io_w_in_15;
  wire  _T_7_io_rdy;
  wire [15:0] _T_7_io_d_out_0;
  wire [15:0] _T_7_io_d_out_1;
  wire [15:0] _T_7_io_d_out_2;
  wire [15:0] _T_7_io_d_out_3;
  wire [15:0] _T_7_io_d_out_4;
  wire [15:0] _T_7_io_d_out_5;
  wire [15:0] _T_7_io_d_out_6;
  wire [15:0] _T_7_io_d_out_7;
  wire [15:0] _T_7_io_d_out_8;
  wire [15:0] _T_7_io_d_out_9;
  wire [15:0] _T_7_io_d_out_10;
  wire [15:0] _T_7_io_d_out_11;
  wire [15:0] _T_7_io_d_out_12;
  wire [15:0] _T_7_io_d_out_13;
  wire [15:0] _T_7_io_d_out_14;
  wire [15:0] _T_7_io_d_out_15;
  wire  _T_7_io_v;
  wire  _T_8_clock;
  wire  _T_8_reset;
  wire [15:0] _T_8_io_d_in;
  wire  _T_8_io_en;
  wire [399:0] _T_8_io_d_out;
  wire  _T_9_clock;
  wire  _T_9_reset;
  wire [399:0] _T_9_io_d_in;
  wire [399:0] _T_9_io_w_in_0;
  wire [399:0] _T_9_io_w_in_1;
  wire [399:0] _T_9_io_w_in_2;
  wire [399:0] _T_9_io_w_in_3;
  wire [399:0] _T_9_io_w_in_4;
  wire [399:0] _T_9_io_w_in_5;
  wire [399:0] _T_9_io_w_in_6;
  wire [399:0] _T_9_io_w_in_7;
  wire [399:0] _T_9_io_w_in_8;
  wire [399:0] _T_9_io_w_in_9;
  wire [399:0] _T_9_io_w_in_10;
  wire [399:0] _T_9_io_w_in_11;
  wire [399:0] _T_9_io_w_in_12;
  wire [399:0] _T_9_io_w_in_13;
  wire [399:0] _T_9_io_w_in_14;
  wire [399:0] _T_9_io_w_in_15;
  wire  _T_9_io_rdy;
  wire [15:0] _T_9_io_d_out_0;
  wire [15:0] _T_9_io_d_out_1;
  wire [15:0] _T_9_io_d_out_2;
  wire [15:0] _T_9_io_d_out_3;
  wire [15:0] _T_9_io_d_out_4;
  wire [15:0] _T_9_io_d_out_5;
  wire [15:0] _T_9_io_d_out_6;
  wire [15:0] _T_9_io_d_out_7;
  wire [15:0] _T_9_io_d_out_8;
  wire [15:0] _T_9_io_d_out_9;
  wire [15:0] _T_9_io_d_out_10;
  wire [15:0] _T_9_io_d_out_11;
  wire [15:0] _T_9_io_d_out_12;
  wire [15:0] _T_9_io_d_out_13;
  wire [15:0] _T_9_io_d_out_14;
  wire [15:0] _T_9_io_d_out_15;
  wire  _T_9_io_v;
  wire  _T_10_clock;
  wire  _T_10_reset;
  wire [15:0] _T_10_io_d_in;
  wire  _T_10_io_en;
  wire [399:0] _T_10_io_d_out;
  wire  _T_11_clock;
  wire  _T_11_reset;
  wire [399:0] _T_11_io_d_in;
  wire [399:0] _T_11_io_w_in_0;
  wire [399:0] _T_11_io_w_in_1;
  wire [399:0] _T_11_io_w_in_2;
  wire [399:0] _T_11_io_w_in_3;
  wire [399:0] _T_11_io_w_in_4;
  wire [399:0] _T_11_io_w_in_5;
  wire [399:0] _T_11_io_w_in_6;
  wire [399:0] _T_11_io_w_in_7;
  wire [399:0] _T_11_io_w_in_8;
  wire [399:0] _T_11_io_w_in_9;
  wire [399:0] _T_11_io_w_in_10;
  wire [399:0] _T_11_io_w_in_11;
  wire [399:0] _T_11_io_w_in_12;
  wire [399:0] _T_11_io_w_in_13;
  wire [399:0] _T_11_io_w_in_14;
  wire [399:0] _T_11_io_w_in_15;
  wire  _T_11_io_rdy;
  wire [15:0] _T_11_io_d_out_0;
  wire [15:0] _T_11_io_d_out_1;
  wire [15:0] _T_11_io_d_out_2;
  wire [15:0] _T_11_io_d_out_3;
  wire [15:0] _T_11_io_d_out_4;
  wire [15:0] _T_11_io_d_out_5;
  wire [15:0] _T_11_io_d_out_6;
  wire [15:0] _T_11_io_d_out_7;
  wire [15:0] _T_11_io_d_out_8;
  wire [15:0] _T_11_io_d_out_9;
  wire [15:0] _T_11_io_d_out_10;
  wire [15:0] _T_11_io_d_out_11;
  wire [15:0] _T_11_io_d_out_12;
  wire [15:0] _T_11_io_d_out_13;
  wire [15:0] _T_11_io_d_out_14;
  wire [15:0] _T_11_io_d_out_15;
  wire  _T_11_io_v;
  reg [15:0] C1_counter;
  reg [31:0] _RAND_0;
  wire  _T_12;
  wire [16:0] _T_13;
  wire [16:0] _GEN_0;
  wire [16:0] _GEN_1;
  wire  _T_14;
  wire  _T_15;
  wire  _T_16;
  wire  _T_17;
  reg [15:0] _T_19;
  reg [31:0] _RAND_1;
  wire [16:0] _T_20;
  wire [16:0] _GEN_3;
  wire [17:0] _T_21;
  wire [17:0] _GEN_4;
  wire [18:0] _T_22;
  wire [18:0] _GEN_5;
  wire [19:0] _T_23;
  wire [19:0] _GEN_6;
  wire [20:0] _T_24;
  wire [21:0] _T_26;
  reg [15:0] _T_27;
  reg [31:0] _RAND_2;
  wire [16:0] _T_28;
  wire [16:0] _GEN_7;
  wire [17:0] _T_29;
  wire [17:0] _GEN_8;
  wire [18:0] _T_30;
  wire [18:0] _GEN_9;
  wire [19:0] _T_31;
  wire [19:0] _GEN_10;
  wire [20:0] _T_32;
  wire [21:0] _T_34;
  reg [15:0] _T_35;
  reg [31:0] _RAND_3;
  wire [16:0] _T_36;
  wire [16:0] _GEN_11;
  wire [17:0] _T_37;
  wire [17:0] _GEN_12;
  wire [18:0] _T_38;
  wire [18:0] _GEN_13;
  wire [19:0] _T_39;
  wire [19:0] _GEN_14;
  wire [20:0] _T_40;
  wire [21:0] _T_42;
  reg [15:0] _T_43;
  reg [31:0] _RAND_4;
  wire [16:0] _T_44;
  wire [16:0] _GEN_15;
  wire [17:0] _T_45;
  wire [17:0] _GEN_16;
  wire [18:0] _T_46;
  wire [18:0] _GEN_17;
  wire [19:0] _T_47;
  wire [19:0] _GEN_18;
  wire [20:0] _T_48;
  wire [21:0] _T_50;
  reg [15:0] _T_51;
  reg [31:0] _RAND_5;
  wire [16:0] _T_52;
  wire [16:0] _GEN_19;
  wire [17:0] _T_53;
  wire [17:0] _GEN_20;
  wire [18:0] _T_54;
  wire [18:0] _GEN_21;
  wire [19:0] _T_55;
  wire [19:0] _GEN_22;
  wire [20:0] _T_56;
  wire [21:0] _T_58;
  reg [15:0] _T_59;
  reg [31:0] _RAND_6;
  wire [16:0] _T_60;
  wire [16:0] _GEN_23;
  wire [17:0] _T_61;
  wire [17:0] _GEN_24;
  wire [18:0] _T_62;
  wire [18:0] _GEN_25;
  wire [19:0] _T_63;
  wire [19:0] _GEN_26;
  wire [20:0] _T_64;
  wire [21:0] _T_66;
  reg [15:0] _T_67;
  reg [31:0] _RAND_7;
  wire [16:0] _T_68;
  wire [16:0] _GEN_27;
  wire [17:0] _T_69;
  wire [17:0] _GEN_28;
  wire [18:0] _T_70;
  wire [18:0] _GEN_29;
  wire [19:0] _T_71;
  wire [19:0] _GEN_30;
  wire [20:0] _T_72;
  wire [21:0] _T_74;
  reg [15:0] _T_75;
  reg [31:0] _RAND_8;
  wire [16:0] _T_76;
  wire [16:0] _GEN_31;
  wire [17:0] _T_77;
  wire [17:0] _GEN_32;
  wire [18:0] _T_78;
  wire [18:0] _GEN_33;
  wire [19:0] _T_79;
  wire [19:0] _GEN_34;
  wire [20:0] _T_80;
  wire [21:0] _T_82;
  reg [15:0] _T_83;
  reg [31:0] _RAND_9;
  wire [16:0] _T_84;
  wire [16:0] _GEN_35;
  wire [17:0] _T_85;
  wire [17:0] _GEN_36;
  wire [18:0] _T_86;
  wire [18:0] _GEN_37;
  wire [19:0] _T_87;
  wire [19:0] _GEN_38;
  wire [20:0] _T_88;
  wire [21:0] _T_90;
  reg [15:0] _T_91;
  reg [31:0] _RAND_10;
  wire [16:0] _T_92;
  wire [16:0] _GEN_39;
  wire [17:0] _T_93;
  wire [17:0] _GEN_40;
  wire [18:0] _T_94;
  wire [18:0] _GEN_41;
  wire [19:0] _T_95;
  wire [19:0] _GEN_42;
  wire [20:0] _T_96;
  wire [21:0] _T_98;
  reg [15:0] _T_99;
  reg [31:0] _RAND_11;
  wire [16:0] _T_100;
  wire [16:0] _GEN_43;
  wire [17:0] _T_101;
  wire [17:0] _GEN_44;
  wire [18:0] _T_102;
  wire [18:0] _GEN_45;
  wire [19:0] _T_103;
  wire [19:0] _GEN_46;
  wire [20:0] _T_104;
  wire [21:0] _T_106;
  reg [15:0] _T_107;
  reg [31:0] _RAND_12;
  wire [16:0] _T_108;
  wire [16:0] _GEN_47;
  wire [17:0] _T_109;
  wire [17:0] _GEN_48;
  wire [18:0] _T_110;
  wire [18:0] _GEN_49;
  wire [19:0] _T_111;
  wire [19:0] _GEN_50;
  wire [20:0] _T_112;
  wire [21:0] _T_114;
  reg [15:0] _T_115;
  reg [31:0] _RAND_13;
  wire [16:0] _T_116;
  wire [16:0] _GEN_51;
  wire [17:0] _T_117;
  wire [17:0] _GEN_52;
  wire [18:0] _T_118;
  wire [18:0] _GEN_53;
  wire [19:0] _T_119;
  wire [19:0] _GEN_54;
  wire [20:0] _T_120;
  wire [21:0] _T_122;
  reg [15:0] _T_123;
  reg [31:0] _RAND_14;
  wire [16:0] _T_124;
  wire [16:0] _GEN_55;
  wire [17:0] _T_125;
  wire [17:0] _GEN_56;
  wire [18:0] _T_126;
  wire [18:0] _GEN_57;
  wire [19:0] _T_127;
  wire [19:0] _GEN_58;
  wire [20:0] _T_128;
  wire [21:0] _T_130;
  reg [15:0] _T_131;
  reg [31:0] _RAND_15;
  wire [16:0] _T_132;
  wire [16:0] _GEN_59;
  wire [17:0] _T_133;
  wire [17:0] _GEN_60;
  wire [18:0] _T_134;
  wire [18:0] _GEN_61;
  wire [19:0] _T_135;
  wire [19:0] _GEN_62;
  wire [20:0] _T_136;
  wire [21:0] _T_138;
  reg [15:0] _T_139;
  reg [31:0] _RAND_16;
  wire [16:0] _T_140;
  wire [16:0] _GEN_63;
  wire [17:0] _T_141;
  wire [17:0] _GEN_64;
  wire [18:0] _T_142;
  wire [18:0] _GEN_65;
  wire [19:0] _T_143;
  wire [19:0] _GEN_66;
  wire [20:0] _T_144;
  wire [21:0] _T_146;
  ShiftRegister _T (
    .clock(_T_clock),
    .reset(_T_reset),
    .io_d_in(_T_io_d_in),
    .io_en(_T_io_en),
    .io_d_out(_T_io_d_out)
  );
  ConvC3 _T_1 (
    .clock(_T_1_clock),
    .reset(_T_1_reset),
    .io_d_in(_T_1_io_d_in),
    .io_w_in_0(_T_1_io_w_in_0),
    .io_w_in_1(_T_1_io_w_in_1),
    .io_w_in_2(_T_1_io_w_in_2),
    .io_w_in_3(_T_1_io_w_in_3),
    .io_w_in_4(_T_1_io_w_in_4),
    .io_w_in_5(_T_1_io_w_in_5),
    .io_w_in_6(_T_1_io_w_in_6),
    .io_w_in_7(_T_1_io_w_in_7),
    .io_w_in_8(_T_1_io_w_in_8),
    .io_w_in_9(_T_1_io_w_in_9),
    .io_w_in_10(_T_1_io_w_in_10),
    .io_w_in_11(_T_1_io_w_in_11),
    .io_w_in_12(_T_1_io_w_in_12),
    .io_w_in_13(_T_1_io_w_in_13),
    .io_w_in_14(_T_1_io_w_in_14),
    .io_w_in_15(_T_1_io_w_in_15),
    .io_rdy(_T_1_io_rdy),
    .io_d_out_0(_T_1_io_d_out_0),
    .io_d_out_1(_T_1_io_d_out_1),
    .io_d_out_2(_T_1_io_d_out_2),
    .io_d_out_3(_T_1_io_d_out_3),
    .io_d_out_4(_T_1_io_d_out_4),
    .io_d_out_5(_T_1_io_d_out_5),
    .io_d_out_6(_T_1_io_d_out_6),
    .io_d_out_7(_T_1_io_d_out_7),
    .io_d_out_8(_T_1_io_d_out_8),
    .io_d_out_9(_T_1_io_d_out_9),
    .io_d_out_10(_T_1_io_d_out_10),
    .io_d_out_11(_T_1_io_d_out_11),
    .io_d_out_12(_T_1_io_d_out_12),
    .io_d_out_13(_T_1_io_d_out_13),
    .io_d_out_14(_T_1_io_d_out_14),
    .io_d_out_15(_T_1_io_d_out_15),
    .io_v(_T_1_io_v)
  );
  ShiftRegister _T_2 (
    .clock(_T_2_clock),
    .reset(_T_2_reset),
    .io_d_in(_T_2_io_d_in),
    .io_en(_T_2_io_en),
    .io_d_out(_T_2_io_d_out)
  );
  ConvC3 _T_3 (
    .clock(_T_3_clock),
    .reset(_T_3_reset),
    .io_d_in(_T_3_io_d_in),
    .io_w_in_0(_T_3_io_w_in_0),
    .io_w_in_1(_T_3_io_w_in_1),
    .io_w_in_2(_T_3_io_w_in_2),
    .io_w_in_3(_T_3_io_w_in_3),
    .io_w_in_4(_T_3_io_w_in_4),
    .io_w_in_5(_T_3_io_w_in_5),
    .io_w_in_6(_T_3_io_w_in_6),
    .io_w_in_7(_T_3_io_w_in_7),
    .io_w_in_8(_T_3_io_w_in_8),
    .io_w_in_9(_T_3_io_w_in_9),
    .io_w_in_10(_T_3_io_w_in_10),
    .io_w_in_11(_T_3_io_w_in_11),
    .io_w_in_12(_T_3_io_w_in_12),
    .io_w_in_13(_T_3_io_w_in_13),
    .io_w_in_14(_T_3_io_w_in_14),
    .io_w_in_15(_T_3_io_w_in_15),
    .io_rdy(_T_3_io_rdy),
    .io_d_out_0(_T_3_io_d_out_0),
    .io_d_out_1(_T_3_io_d_out_1),
    .io_d_out_2(_T_3_io_d_out_2),
    .io_d_out_3(_T_3_io_d_out_3),
    .io_d_out_4(_T_3_io_d_out_4),
    .io_d_out_5(_T_3_io_d_out_5),
    .io_d_out_6(_T_3_io_d_out_6),
    .io_d_out_7(_T_3_io_d_out_7),
    .io_d_out_8(_T_3_io_d_out_8),
    .io_d_out_9(_T_3_io_d_out_9),
    .io_d_out_10(_T_3_io_d_out_10),
    .io_d_out_11(_T_3_io_d_out_11),
    .io_d_out_12(_T_3_io_d_out_12),
    .io_d_out_13(_T_3_io_d_out_13),
    .io_d_out_14(_T_3_io_d_out_14),
    .io_d_out_15(_T_3_io_d_out_15),
    .io_v(_T_3_io_v)
  );
  ShiftRegister _T_4 (
    .clock(_T_4_clock),
    .reset(_T_4_reset),
    .io_d_in(_T_4_io_d_in),
    .io_en(_T_4_io_en),
    .io_d_out(_T_4_io_d_out)
  );
  ConvC3 _T_5 (
    .clock(_T_5_clock),
    .reset(_T_5_reset),
    .io_d_in(_T_5_io_d_in),
    .io_w_in_0(_T_5_io_w_in_0),
    .io_w_in_1(_T_5_io_w_in_1),
    .io_w_in_2(_T_5_io_w_in_2),
    .io_w_in_3(_T_5_io_w_in_3),
    .io_w_in_4(_T_5_io_w_in_4),
    .io_w_in_5(_T_5_io_w_in_5),
    .io_w_in_6(_T_5_io_w_in_6),
    .io_w_in_7(_T_5_io_w_in_7),
    .io_w_in_8(_T_5_io_w_in_8),
    .io_w_in_9(_T_5_io_w_in_9),
    .io_w_in_10(_T_5_io_w_in_10),
    .io_w_in_11(_T_5_io_w_in_11),
    .io_w_in_12(_T_5_io_w_in_12),
    .io_w_in_13(_T_5_io_w_in_13),
    .io_w_in_14(_T_5_io_w_in_14),
    .io_w_in_15(_T_5_io_w_in_15),
    .io_rdy(_T_5_io_rdy),
    .io_d_out_0(_T_5_io_d_out_0),
    .io_d_out_1(_T_5_io_d_out_1),
    .io_d_out_2(_T_5_io_d_out_2),
    .io_d_out_3(_T_5_io_d_out_3),
    .io_d_out_4(_T_5_io_d_out_4),
    .io_d_out_5(_T_5_io_d_out_5),
    .io_d_out_6(_T_5_io_d_out_6),
    .io_d_out_7(_T_5_io_d_out_7),
    .io_d_out_8(_T_5_io_d_out_8),
    .io_d_out_9(_T_5_io_d_out_9),
    .io_d_out_10(_T_5_io_d_out_10),
    .io_d_out_11(_T_5_io_d_out_11),
    .io_d_out_12(_T_5_io_d_out_12),
    .io_d_out_13(_T_5_io_d_out_13),
    .io_d_out_14(_T_5_io_d_out_14),
    .io_d_out_15(_T_5_io_d_out_15),
    .io_v(_T_5_io_v)
  );
  ShiftRegister _T_6 (
    .clock(_T_6_clock),
    .reset(_T_6_reset),
    .io_d_in(_T_6_io_d_in),
    .io_en(_T_6_io_en),
    .io_d_out(_T_6_io_d_out)
  );
  ConvC3 _T_7 (
    .clock(_T_7_clock),
    .reset(_T_7_reset),
    .io_d_in(_T_7_io_d_in),
    .io_w_in_0(_T_7_io_w_in_0),
    .io_w_in_1(_T_7_io_w_in_1),
    .io_w_in_2(_T_7_io_w_in_2),
    .io_w_in_3(_T_7_io_w_in_3),
    .io_w_in_4(_T_7_io_w_in_4),
    .io_w_in_5(_T_7_io_w_in_5),
    .io_w_in_6(_T_7_io_w_in_6),
    .io_w_in_7(_T_7_io_w_in_7),
    .io_w_in_8(_T_7_io_w_in_8),
    .io_w_in_9(_T_7_io_w_in_9),
    .io_w_in_10(_T_7_io_w_in_10),
    .io_w_in_11(_T_7_io_w_in_11),
    .io_w_in_12(_T_7_io_w_in_12),
    .io_w_in_13(_T_7_io_w_in_13),
    .io_w_in_14(_T_7_io_w_in_14),
    .io_w_in_15(_T_7_io_w_in_15),
    .io_rdy(_T_7_io_rdy),
    .io_d_out_0(_T_7_io_d_out_0),
    .io_d_out_1(_T_7_io_d_out_1),
    .io_d_out_2(_T_7_io_d_out_2),
    .io_d_out_3(_T_7_io_d_out_3),
    .io_d_out_4(_T_7_io_d_out_4),
    .io_d_out_5(_T_7_io_d_out_5),
    .io_d_out_6(_T_7_io_d_out_6),
    .io_d_out_7(_T_7_io_d_out_7),
    .io_d_out_8(_T_7_io_d_out_8),
    .io_d_out_9(_T_7_io_d_out_9),
    .io_d_out_10(_T_7_io_d_out_10),
    .io_d_out_11(_T_7_io_d_out_11),
    .io_d_out_12(_T_7_io_d_out_12),
    .io_d_out_13(_T_7_io_d_out_13),
    .io_d_out_14(_T_7_io_d_out_14),
    .io_d_out_15(_T_7_io_d_out_15),
    .io_v(_T_7_io_v)
  );
  ShiftRegister _T_8 (
    .clock(_T_8_clock),
    .reset(_T_8_reset),
    .io_d_in(_T_8_io_d_in),
    .io_en(_T_8_io_en),
    .io_d_out(_T_8_io_d_out)
  );
  ConvC3 _T_9 (
    .clock(_T_9_clock),
    .reset(_T_9_reset),
    .io_d_in(_T_9_io_d_in),
    .io_w_in_0(_T_9_io_w_in_0),
    .io_w_in_1(_T_9_io_w_in_1),
    .io_w_in_2(_T_9_io_w_in_2),
    .io_w_in_3(_T_9_io_w_in_3),
    .io_w_in_4(_T_9_io_w_in_4),
    .io_w_in_5(_T_9_io_w_in_5),
    .io_w_in_6(_T_9_io_w_in_6),
    .io_w_in_7(_T_9_io_w_in_7),
    .io_w_in_8(_T_9_io_w_in_8),
    .io_w_in_9(_T_9_io_w_in_9),
    .io_w_in_10(_T_9_io_w_in_10),
    .io_w_in_11(_T_9_io_w_in_11),
    .io_w_in_12(_T_9_io_w_in_12),
    .io_w_in_13(_T_9_io_w_in_13),
    .io_w_in_14(_T_9_io_w_in_14),
    .io_w_in_15(_T_9_io_w_in_15),
    .io_rdy(_T_9_io_rdy),
    .io_d_out_0(_T_9_io_d_out_0),
    .io_d_out_1(_T_9_io_d_out_1),
    .io_d_out_2(_T_9_io_d_out_2),
    .io_d_out_3(_T_9_io_d_out_3),
    .io_d_out_4(_T_9_io_d_out_4),
    .io_d_out_5(_T_9_io_d_out_5),
    .io_d_out_6(_T_9_io_d_out_6),
    .io_d_out_7(_T_9_io_d_out_7),
    .io_d_out_8(_T_9_io_d_out_8),
    .io_d_out_9(_T_9_io_d_out_9),
    .io_d_out_10(_T_9_io_d_out_10),
    .io_d_out_11(_T_9_io_d_out_11),
    .io_d_out_12(_T_9_io_d_out_12),
    .io_d_out_13(_T_9_io_d_out_13),
    .io_d_out_14(_T_9_io_d_out_14),
    .io_d_out_15(_T_9_io_d_out_15),
    .io_v(_T_9_io_v)
  );
  ShiftRegister _T_10 (
    .clock(_T_10_clock),
    .reset(_T_10_reset),
    .io_d_in(_T_10_io_d_in),
    .io_en(_T_10_io_en),
    .io_d_out(_T_10_io_d_out)
  );
  ConvC3 _T_11 (
    .clock(_T_11_clock),
    .reset(_T_11_reset),
    .io_d_in(_T_11_io_d_in),
    .io_w_in_0(_T_11_io_w_in_0),
    .io_w_in_1(_T_11_io_w_in_1),
    .io_w_in_2(_T_11_io_w_in_2),
    .io_w_in_3(_T_11_io_w_in_3),
    .io_w_in_4(_T_11_io_w_in_4),
    .io_w_in_5(_T_11_io_w_in_5),
    .io_w_in_6(_T_11_io_w_in_6),
    .io_w_in_7(_T_11_io_w_in_7),
    .io_w_in_8(_T_11_io_w_in_8),
    .io_w_in_9(_T_11_io_w_in_9),
    .io_w_in_10(_T_11_io_w_in_10),
    .io_w_in_11(_T_11_io_w_in_11),
    .io_w_in_12(_T_11_io_w_in_12),
    .io_w_in_13(_T_11_io_w_in_13),
    .io_w_in_14(_T_11_io_w_in_14),
    .io_w_in_15(_T_11_io_w_in_15),
    .io_rdy(_T_11_io_rdy),
    .io_d_out_0(_T_11_io_d_out_0),
    .io_d_out_1(_T_11_io_d_out_1),
    .io_d_out_2(_T_11_io_d_out_2),
    .io_d_out_3(_T_11_io_d_out_3),
    .io_d_out_4(_T_11_io_d_out_4),
    .io_d_out_5(_T_11_io_d_out_5),
    .io_d_out_6(_T_11_io_d_out_6),
    .io_d_out_7(_T_11_io_d_out_7),
    .io_d_out_8(_T_11_io_d_out_8),
    .io_d_out_9(_T_11_io_d_out_9),
    .io_d_out_10(_T_11_io_d_out_10),
    .io_d_out_11(_T_11_io_d_out_11),
    .io_d_out_12(_T_11_io_d_out_12),
    .io_d_out_13(_T_11_io_d_out_13),
    .io_d_out_14(_T_11_io_d_out_14),
    .io_d_out_15(_T_11_io_d_out_15),
    .io_v(_T_11_io_v)
  );
  assign _T_12 = C1_counter == 16'h19;
  assign _T_13 = C1_counter + 16'h1;
  assign _GEN_0 = io_rdy ? _T_13 : {{1'd0}, C1_counter};
  assign _GEN_1 = _T_12 ? 17'h0 : _GEN_0;
  assign _T_14 = _T_1_io_v & _T_3_io_v;
  assign _T_15 = _T_14 & _T_5_io_v;
  assign _T_16 = _T_15 & _T_7_io_v;
  assign _T_17 = _T_16 & _T_9_io_v;
  assign _T_20 = _T_1_io_d_out_0 + _T_3_io_d_out_0;
  assign _GEN_3 = {{1'd0}, _T_5_io_d_out_0};
  assign _T_21 = _T_20 + _GEN_3;
  assign _GEN_4 = {{2'd0}, _T_7_io_d_out_0};
  assign _T_22 = _T_21 + _GEN_4;
  assign _GEN_5 = {{3'd0}, _T_9_io_d_out_0};
  assign _T_23 = _T_22 + _GEN_5;
  assign _GEN_6 = {{4'd0}, _T_11_io_d_out_0};
  assign _T_24 = _T_23 + _GEN_6;
  assign _T_26 = _T_24 + 21'h1;
  assign _T_28 = _T_1_io_d_out_1 + _T_3_io_d_out_1;
  assign _GEN_7 = {{1'd0}, _T_5_io_d_out_1};
  assign _T_29 = _T_28 + _GEN_7;
  assign _GEN_8 = {{2'd0}, _T_7_io_d_out_1};
  assign _T_30 = _T_29 + _GEN_8;
  assign _GEN_9 = {{3'd0}, _T_9_io_d_out_1};
  assign _T_31 = _T_30 + _GEN_9;
  assign _GEN_10 = {{4'd0}, _T_11_io_d_out_1};
  assign _T_32 = _T_31 + _GEN_10;
  assign _T_34 = {{1'd0}, _T_32};
  assign _T_36 = _T_1_io_d_out_2 + _T_3_io_d_out_2;
  assign _GEN_11 = {{1'd0}, _T_5_io_d_out_2};
  assign _T_37 = _T_36 + _GEN_11;
  assign _GEN_12 = {{2'd0}, _T_7_io_d_out_2};
  assign _T_38 = _T_37 + _GEN_12;
  assign _GEN_13 = {{3'd0}, _T_9_io_d_out_2};
  assign _T_39 = _T_38 + _GEN_13;
  assign _GEN_14 = {{4'd0}, _T_11_io_d_out_2};
  assign _T_40 = _T_39 + _GEN_14;
  assign _T_42 = {{1'd0}, _T_40};
  assign _T_44 = _T_1_io_d_out_3 + _T_3_io_d_out_3;
  assign _GEN_15 = {{1'd0}, _T_5_io_d_out_3};
  assign _T_45 = _T_44 + _GEN_15;
  assign _GEN_16 = {{2'd0}, _T_7_io_d_out_3};
  assign _T_46 = _T_45 + _GEN_16;
  assign _GEN_17 = {{3'd0}, _T_9_io_d_out_3};
  assign _T_47 = _T_46 + _GEN_17;
  assign _GEN_18 = {{4'd0}, _T_11_io_d_out_3};
  assign _T_48 = _T_47 + _GEN_18;
  assign _T_50 = {{1'd0}, _T_48};
  assign _T_52 = _T_1_io_d_out_4 + _T_3_io_d_out_4;
  assign _GEN_19 = {{1'd0}, _T_5_io_d_out_4};
  assign _T_53 = _T_52 + _GEN_19;
  assign _GEN_20 = {{2'd0}, _T_7_io_d_out_4};
  assign _T_54 = _T_53 + _GEN_20;
  assign _GEN_21 = {{3'd0}, _T_9_io_d_out_4};
  assign _T_55 = _T_54 + _GEN_21;
  assign _GEN_22 = {{4'd0}, _T_11_io_d_out_4};
  assign _T_56 = _T_55 + _GEN_22;
  assign _T_58 = {{1'd0}, _T_56};
  assign _T_60 = _T_1_io_d_out_5 + _T_3_io_d_out_5;
  assign _GEN_23 = {{1'd0}, _T_5_io_d_out_5};
  assign _T_61 = _T_60 + _GEN_23;
  assign _GEN_24 = {{2'd0}, _T_7_io_d_out_5};
  assign _T_62 = _T_61 + _GEN_24;
  assign _GEN_25 = {{3'd0}, _T_9_io_d_out_5};
  assign _T_63 = _T_62 + _GEN_25;
  assign _GEN_26 = {{4'd0}, _T_11_io_d_out_5};
  assign _T_64 = _T_63 + _GEN_26;
  assign _T_66 = {{1'd0}, _T_64};
  assign _T_68 = _T_1_io_d_out_6 + _T_3_io_d_out_6;
  assign _GEN_27 = {{1'd0}, _T_5_io_d_out_6};
  assign _T_69 = _T_68 + _GEN_27;
  assign _GEN_28 = {{2'd0}, _T_7_io_d_out_6};
  assign _T_70 = _T_69 + _GEN_28;
  assign _GEN_29 = {{3'd0}, _T_9_io_d_out_6};
  assign _T_71 = _T_70 + _GEN_29;
  assign _GEN_30 = {{4'd0}, _T_11_io_d_out_6};
  assign _T_72 = _T_71 + _GEN_30;
  assign _T_74 = {{1'd0}, _T_72};
  assign _T_76 = _T_1_io_d_out_7 + _T_3_io_d_out_7;
  assign _GEN_31 = {{1'd0}, _T_5_io_d_out_7};
  assign _T_77 = _T_76 + _GEN_31;
  assign _GEN_32 = {{2'd0}, _T_7_io_d_out_7};
  assign _T_78 = _T_77 + _GEN_32;
  assign _GEN_33 = {{3'd0}, _T_9_io_d_out_7};
  assign _T_79 = _T_78 + _GEN_33;
  assign _GEN_34 = {{4'd0}, _T_11_io_d_out_7};
  assign _T_80 = _T_79 + _GEN_34;
  assign _T_82 = {{1'd0}, _T_80};
  assign _T_84 = _T_1_io_d_out_8 + _T_3_io_d_out_8;
  assign _GEN_35 = {{1'd0}, _T_5_io_d_out_8};
  assign _T_85 = _T_84 + _GEN_35;
  assign _GEN_36 = {{2'd0}, _T_7_io_d_out_8};
  assign _T_86 = _T_85 + _GEN_36;
  assign _GEN_37 = {{3'd0}, _T_9_io_d_out_8};
  assign _T_87 = _T_86 + _GEN_37;
  assign _GEN_38 = {{4'd0}, _T_11_io_d_out_8};
  assign _T_88 = _T_87 + _GEN_38;
  assign _T_90 = {{1'd0}, _T_88};
  assign _T_92 = _T_1_io_d_out_9 + _T_3_io_d_out_9;
  assign _GEN_39 = {{1'd0}, _T_5_io_d_out_9};
  assign _T_93 = _T_92 + _GEN_39;
  assign _GEN_40 = {{2'd0}, _T_7_io_d_out_9};
  assign _T_94 = _T_93 + _GEN_40;
  assign _GEN_41 = {{3'd0}, _T_9_io_d_out_9};
  assign _T_95 = _T_94 + _GEN_41;
  assign _GEN_42 = {{4'd0}, _T_11_io_d_out_9};
  assign _T_96 = _T_95 + _GEN_42;
  assign _T_98 = {{1'd0}, _T_96};
  assign _T_100 = _T_1_io_d_out_10 + _T_3_io_d_out_10;
  assign _GEN_43 = {{1'd0}, _T_5_io_d_out_10};
  assign _T_101 = _T_100 + _GEN_43;
  assign _GEN_44 = {{2'd0}, _T_7_io_d_out_10};
  assign _T_102 = _T_101 + _GEN_44;
  assign _GEN_45 = {{3'd0}, _T_9_io_d_out_10};
  assign _T_103 = _T_102 + _GEN_45;
  assign _GEN_46 = {{4'd0}, _T_11_io_d_out_10};
  assign _T_104 = _T_103 + _GEN_46;
  assign _T_106 = {{1'd0}, _T_104};
  assign _T_108 = _T_1_io_d_out_11 + _T_3_io_d_out_11;
  assign _GEN_47 = {{1'd0}, _T_5_io_d_out_11};
  assign _T_109 = _T_108 + _GEN_47;
  assign _GEN_48 = {{2'd0}, _T_7_io_d_out_11};
  assign _T_110 = _T_109 + _GEN_48;
  assign _GEN_49 = {{3'd0}, _T_9_io_d_out_11};
  assign _T_111 = _T_110 + _GEN_49;
  assign _GEN_50 = {{4'd0}, _T_11_io_d_out_11};
  assign _T_112 = _T_111 + _GEN_50;
  assign _T_114 = {{1'd0}, _T_112};
  assign _T_116 = _T_1_io_d_out_12 + _T_3_io_d_out_12;
  assign _GEN_51 = {{1'd0}, _T_5_io_d_out_12};
  assign _T_117 = _T_116 + _GEN_51;
  assign _GEN_52 = {{2'd0}, _T_7_io_d_out_12};
  assign _T_118 = _T_117 + _GEN_52;
  assign _GEN_53 = {{3'd0}, _T_9_io_d_out_12};
  assign _T_119 = _T_118 + _GEN_53;
  assign _GEN_54 = {{4'd0}, _T_11_io_d_out_12};
  assign _T_120 = _T_119 + _GEN_54;
  assign _T_122 = {{1'd0}, _T_120};
  assign _T_124 = _T_1_io_d_out_13 + _T_3_io_d_out_13;
  assign _GEN_55 = {{1'd0}, _T_5_io_d_out_13};
  assign _T_125 = _T_124 + _GEN_55;
  assign _GEN_56 = {{2'd0}, _T_7_io_d_out_13};
  assign _T_126 = _T_125 + _GEN_56;
  assign _GEN_57 = {{3'd0}, _T_9_io_d_out_13};
  assign _T_127 = _T_126 + _GEN_57;
  assign _GEN_58 = {{4'd0}, _T_11_io_d_out_13};
  assign _T_128 = _T_127 + _GEN_58;
  assign _T_130 = {{1'd0}, _T_128};
  assign _T_132 = _T_1_io_d_out_14 + _T_3_io_d_out_14;
  assign _GEN_59 = {{1'd0}, _T_5_io_d_out_14};
  assign _T_133 = _T_132 + _GEN_59;
  assign _GEN_60 = {{2'd0}, _T_7_io_d_out_14};
  assign _T_134 = _T_133 + _GEN_60;
  assign _GEN_61 = {{3'd0}, _T_9_io_d_out_14};
  assign _T_135 = _T_134 + _GEN_61;
  assign _GEN_62 = {{4'd0}, _T_11_io_d_out_14};
  assign _T_136 = _T_135 + _GEN_62;
  assign _T_138 = {{1'd0}, _T_136};
  assign _T_140 = _T_1_io_d_out_15 + _T_3_io_d_out_15;
  assign _GEN_63 = {{1'd0}, _T_5_io_d_out_15};
  assign _T_141 = _T_140 + _GEN_63;
  assign _GEN_64 = {{2'd0}, _T_7_io_d_out_15};
  assign _T_142 = _T_141 + _GEN_64;
  assign _GEN_65 = {{3'd0}, _T_9_io_d_out_15};
  assign _T_143 = _T_142 + _GEN_65;
  assign _GEN_66 = {{4'd0}, _T_11_io_d_out_15};
  assign _T_144 = _T_143 + _GEN_66;
  assign _T_146 = {{1'd0}, _T_144};
  assign io_c3_v = _T_17 & _T_11_io_v;
  assign io_d_out_0 = _T_19;
  assign io_d_out_1 = _T_27;
  assign io_d_out_2 = _T_35;
  assign io_d_out_3 = _T_43;
  assign io_d_out_4 = _T_51;
  assign io_d_out_5 = _T_59;
  assign io_d_out_6 = _T_67;
  assign io_d_out_7 = _T_75;
  assign io_d_out_8 = _T_83;
  assign io_d_out_9 = _T_91;
  assign io_d_out_10 = _T_99;
  assign io_d_out_11 = _T_107;
  assign io_d_out_12 = _T_115;
  assign io_d_out_13 = _T_123;
  assign io_d_out_14 = _T_131;
  assign io_d_out_15 = _T_139;
  assign _T_clock = clock;
  assign _T_reset = reset;
  assign _T_io_d_in = io_d_in_0;
  assign _T_io_en = io_rdy;
  assign _T_1_clock = clock;
  assign _T_1_reset = reset;
  assign _T_1_io_d_in = _T_io_d_out;
  assign _T_1_io_w_in_0 = 400'h0;
  assign _T_1_io_w_in_1 = 400'h0;
  assign _T_1_io_w_in_2 = 400'h0;
  assign _T_1_io_w_in_3 = 400'h0;
  assign _T_1_io_w_in_4 = 400'h0;
  assign _T_1_io_w_in_5 = 400'h0;
  assign _T_1_io_w_in_6 = 400'h0;
  assign _T_1_io_w_in_7 = 400'h0;
  assign _T_1_io_w_in_8 = 400'h0;
  assign _T_1_io_w_in_9 = 400'h0;
  assign _T_1_io_w_in_10 = 400'h0;
  assign _T_1_io_w_in_11 = 400'h0;
  assign _T_1_io_w_in_12 = 400'h0;
  assign _T_1_io_w_in_13 = 400'h0;
  assign _T_1_io_w_in_14 = 400'h0;
  assign _T_1_io_w_in_15 = 400'h0;
  assign _T_1_io_rdy = C1_counter == 16'h19;
  assign _T_2_clock = clock;
  assign _T_2_reset = reset;
  assign _T_2_io_d_in = io_d_in_1;
  assign _T_2_io_en = io_rdy;
  assign _T_3_clock = clock;
  assign _T_3_reset = reset;
  assign _T_3_io_d_in = _T_2_io_d_out;
  assign _T_3_io_w_in_0 = 400'h1;
  assign _T_3_io_w_in_1 = 400'h1;
  assign _T_3_io_w_in_2 = 400'h1;
  assign _T_3_io_w_in_3 = 400'h1;
  assign _T_3_io_w_in_4 = 400'h1;
  assign _T_3_io_w_in_5 = 400'h1;
  assign _T_3_io_w_in_6 = 400'h1;
  assign _T_3_io_w_in_7 = 400'h1;
  assign _T_3_io_w_in_8 = 400'h1;
  assign _T_3_io_w_in_9 = 400'h1;
  assign _T_3_io_w_in_10 = 400'h1;
  assign _T_3_io_w_in_11 = 400'h1;
  assign _T_3_io_w_in_12 = 400'h1;
  assign _T_3_io_w_in_13 = 400'h1;
  assign _T_3_io_w_in_14 = 400'h1;
  assign _T_3_io_w_in_15 = 400'h1;
  assign _T_3_io_rdy = C1_counter == 16'h19;
  assign _T_4_clock = clock;
  assign _T_4_reset = reset;
  assign _T_4_io_d_in = io_d_in_2;
  assign _T_4_io_en = io_rdy;
  assign _T_5_clock = clock;
  assign _T_5_reset = reset;
  assign _T_5_io_d_in = _T_4_io_d_out;
  assign _T_5_io_w_in_0 = 400'h2;
  assign _T_5_io_w_in_1 = 400'h2;
  assign _T_5_io_w_in_2 = 400'h2;
  assign _T_5_io_w_in_3 = 400'h2;
  assign _T_5_io_w_in_4 = 400'h2;
  assign _T_5_io_w_in_5 = 400'h2;
  assign _T_5_io_w_in_6 = 400'h2;
  assign _T_5_io_w_in_7 = 400'h2;
  assign _T_5_io_w_in_8 = 400'h2;
  assign _T_5_io_w_in_9 = 400'h2;
  assign _T_5_io_w_in_10 = 400'h2;
  assign _T_5_io_w_in_11 = 400'h2;
  assign _T_5_io_w_in_12 = 400'h2;
  assign _T_5_io_w_in_13 = 400'h2;
  assign _T_5_io_w_in_14 = 400'h2;
  assign _T_5_io_w_in_15 = 400'h2;
  assign _T_5_io_rdy = C1_counter == 16'h19;
  assign _T_6_clock = clock;
  assign _T_6_reset = reset;
  assign _T_6_io_d_in = io_d_in_3;
  assign _T_6_io_en = io_rdy;
  assign _T_7_clock = clock;
  assign _T_7_reset = reset;
  assign _T_7_io_d_in = _T_6_io_d_out;
  assign _T_7_io_w_in_0 = 400'h3;
  assign _T_7_io_w_in_1 = 400'h3;
  assign _T_7_io_w_in_2 = 400'h3;
  assign _T_7_io_w_in_3 = 400'h3;
  assign _T_7_io_w_in_4 = 400'h3;
  assign _T_7_io_w_in_5 = 400'h3;
  assign _T_7_io_w_in_6 = 400'h3;
  assign _T_7_io_w_in_7 = 400'h3;
  assign _T_7_io_w_in_8 = 400'h3;
  assign _T_7_io_w_in_9 = 400'h3;
  assign _T_7_io_w_in_10 = 400'h3;
  assign _T_7_io_w_in_11 = 400'h3;
  assign _T_7_io_w_in_12 = 400'h3;
  assign _T_7_io_w_in_13 = 400'h3;
  assign _T_7_io_w_in_14 = 400'h3;
  assign _T_7_io_w_in_15 = 400'h3;
  assign _T_7_io_rdy = C1_counter == 16'h19;
  assign _T_8_clock = clock;
  assign _T_8_reset = reset;
  assign _T_8_io_d_in = io_d_in_4;
  assign _T_8_io_en = io_rdy;
  assign _T_9_clock = clock;
  assign _T_9_reset = reset;
  assign _T_9_io_d_in = _T_8_io_d_out;
  assign _T_9_io_w_in_0 = 400'h4;
  assign _T_9_io_w_in_1 = 400'h4;
  assign _T_9_io_w_in_2 = 400'h4;
  assign _T_9_io_w_in_3 = 400'h4;
  assign _T_9_io_w_in_4 = 400'h4;
  assign _T_9_io_w_in_5 = 400'h4;
  assign _T_9_io_w_in_6 = 400'h4;
  assign _T_9_io_w_in_7 = 400'h4;
  assign _T_9_io_w_in_8 = 400'h4;
  assign _T_9_io_w_in_9 = 400'h4;
  assign _T_9_io_w_in_10 = 400'h4;
  assign _T_9_io_w_in_11 = 400'h4;
  assign _T_9_io_w_in_12 = 400'h4;
  assign _T_9_io_w_in_13 = 400'h4;
  assign _T_9_io_w_in_14 = 400'h4;
  assign _T_9_io_w_in_15 = 400'h4;
  assign _T_9_io_rdy = C1_counter == 16'h19;
  assign _T_10_clock = clock;
  assign _T_10_reset = reset;
  assign _T_10_io_d_in = io_d_in_5;
  assign _T_10_io_en = io_rdy;
  assign _T_11_clock = clock;
  assign _T_11_reset = reset;
  assign _T_11_io_d_in = _T_10_io_d_out;
  assign _T_11_io_w_in_0 = 400'h5;
  assign _T_11_io_w_in_1 = 400'h5;
  assign _T_11_io_w_in_2 = 400'h5;
  assign _T_11_io_w_in_3 = 400'h5;
  assign _T_11_io_w_in_4 = 400'h5;
  assign _T_11_io_w_in_5 = 400'h5;
  assign _T_11_io_w_in_6 = 400'h5;
  assign _T_11_io_w_in_7 = 400'h5;
  assign _T_11_io_w_in_8 = 400'h5;
  assign _T_11_io_w_in_9 = 400'h5;
  assign _T_11_io_w_in_10 = 400'h5;
  assign _T_11_io_w_in_11 = 400'h5;
  assign _T_11_io_w_in_12 = 400'h5;
  assign _T_11_io_w_in_13 = 400'h5;
  assign _T_11_io_w_in_14 = 400'h5;
  assign _T_11_io_w_in_15 = 400'h5;
  assign _T_11_io_rdy = C1_counter == 16'h19;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  C1_counter = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_19 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_27 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_35 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_43 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_51 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_59 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_67 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_75 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_83 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_91 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_99 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_107 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_115 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_123 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_131 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_139 = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      C1_counter <= 16'h0;
    end else begin
      C1_counter <= _GEN_1[15:0];
    end
    if (reset) begin
      _T_19 <= 16'h0;
    end else begin
      _T_19 <= _T_26[15:0];
    end
    if (reset) begin
      _T_27 <= 16'h0;
    end else begin
      _T_27 <= _T_34[15:0];
    end
    if (reset) begin
      _T_35 <= 16'h0;
    end else begin
      _T_35 <= _T_42[15:0];
    end
    if (reset) begin
      _T_43 <= 16'h0;
    end else begin
      _T_43 <= _T_50[15:0];
    end
    if (reset) begin
      _T_51 <= 16'h0;
    end else begin
      _T_51 <= _T_58[15:0];
    end
    if (reset) begin
      _T_59 <= 16'h0;
    end else begin
      _T_59 <= _T_66[15:0];
    end
    if (reset) begin
      _T_67 <= 16'h0;
    end else begin
      _T_67 <= _T_74[15:0];
    end
    if (reset) begin
      _T_75 <= 16'h0;
    end else begin
      _T_75 <= _T_82[15:0];
    end
    if (reset) begin
      _T_83 <= 16'h0;
    end else begin
      _T_83 <= _T_90[15:0];
    end
    if (reset) begin
      _T_91 <= 16'h0;
    end else begin
      _T_91 <= _T_98[15:0];
    end
    if (reset) begin
      _T_99 <= 16'h0;
    end else begin
      _T_99 <= _T_106[15:0];
    end
    if (reset) begin
      _T_107 <= 16'h0;
    end else begin
      _T_107 <= _T_114[15:0];
    end
    if (reset) begin
      _T_115 <= 16'h0;
    end else begin
      _T_115 <= _T_122[15:0];
    end
    if (reset) begin
      _T_123 <= 16'h0;
    end else begin
      _T_123 <= _T_130[15:0];
    end
    if (reset) begin
      _T_131 <= 16'h0;
    end else begin
      _T_131 <= _T_138[15:0];
    end
    if (reset) begin
      _T_139 <= 16'h0;
    end else begin
      _T_139 <= _T_146[15:0];
    end
  end
endmodule
module C2MaxPool(
  input         clock,
  input         reset,
  input  [15:0] io_d_in_0,
  input  [15:0] io_d_in_1,
  input  [15:0] io_d_in_2,
  input  [15:0] io_d_in_3,
  input  [15:0] io_d_in_4,
  input  [15:0] io_d_in_5,
  input  [15:0] io_d_in_6,
  input  [15:0] io_d_in_7,
  input  [15:0] io_d_in_8,
  input  [15:0] io_d_in_9,
  input  [15:0] io_d_in_10,
  input  [15:0] io_d_in_11,
  input  [15:0] io_d_in_12,
  input  [15:0] io_d_in_13,
  input  [15:0] io_d_in_14,
  input  [15:0] io_d_in_15,
  input         io_rdy,
  output [15:0] io_d_out_0,
  output [15:0] io_d_out_1,
  output [15:0] io_d_out_2,
  output [15:0] io_d_out_3,
  output [15:0] io_d_out_4,
  output [15:0] io_d_out_5,
  output [15:0] io_d_out_6,
  output [15:0] io_d_out_7,
  output [15:0] io_d_out_8,
  output [15:0] io_d_out_9,
  output [15:0] io_d_out_10,
  output [15:0] io_d_out_11,
  output [15:0] io_d_out_12,
  output [15:0] io_d_out_13,
  output [15:0] io_d_out_14,
  output [15:0] io_d_out_15,
  output        io_pool_v
);
  wire  _T_clock;
  wire  _T_reset;
  wire [15:0] _T_io_d_in;
  wire  _T_io_rdy;
  wire [15:0] _T_io_d_out;
  wire  _T_io_v;
  wire  _T_1_clock;
  wire  _T_1_reset;
  wire [15:0] _T_1_io_d_in;
  wire  _T_1_io_rdy;
  wire [15:0] _T_1_io_d_out;
  wire  _T_1_io_v;
  wire  _T_2_clock;
  wire  _T_2_reset;
  wire [15:0] _T_2_io_d_in;
  wire  _T_2_io_rdy;
  wire [15:0] _T_2_io_d_out;
  wire  _T_2_io_v;
  wire  _T_3_clock;
  wire  _T_3_reset;
  wire [15:0] _T_3_io_d_in;
  wire  _T_3_io_rdy;
  wire [15:0] _T_3_io_d_out;
  wire  _T_3_io_v;
  wire  _T_4_clock;
  wire  _T_4_reset;
  wire [15:0] _T_4_io_d_in;
  wire  _T_4_io_rdy;
  wire [15:0] _T_4_io_d_out;
  wire  _T_4_io_v;
  wire  _T_5_clock;
  wire  _T_5_reset;
  wire [15:0] _T_5_io_d_in;
  wire  _T_5_io_rdy;
  wire [15:0] _T_5_io_d_out;
  wire  _T_5_io_v;
  wire  _T_6_clock;
  wire  _T_6_reset;
  wire [15:0] _T_6_io_d_in;
  wire  _T_6_io_rdy;
  wire [15:0] _T_6_io_d_out;
  wire  _T_6_io_v;
  wire  _T_7_clock;
  wire  _T_7_reset;
  wire [15:0] _T_7_io_d_in;
  wire  _T_7_io_rdy;
  wire [15:0] _T_7_io_d_out;
  wire  _T_7_io_v;
  wire  _T_8_clock;
  wire  _T_8_reset;
  wire [15:0] _T_8_io_d_in;
  wire  _T_8_io_rdy;
  wire [15:0] _T_8_io_d_out;
  wire  _T_8_io_v;
  wire  _T_9_clock;
  wire  _T_9_reset;
  wire [15:0] _T_9_io_d_in;
  wire  _T_9_io_rdy;
  wire [15:0] _T_9_io_d_out;
  wire  _T_9_io_v;
  wire  _T_10_clock;
  wire  _T_10_reset;
  wire [15:0] _T_10_io_d_in;
  wire  _T_10_io_rdy;
  wire [15:0] _T_10_io_d_out;
  wire  _T_10_io_v;
  wire  _T_11_clock;
  wire  _T_11_reset;
  wire [15:0] _T_11_io_d_in;
  wire  _T_11_io_rdy;
  wire [15:0] _T_11_io_d_out;
  wire  _T_11_io_v;
  wire  _T_12_clock;
  wire  _T_12_reset;
  wire [15:0] _T_12_io_d_in;
  wire  _T_12_io_rdy;
  wire [15:0] _T_12_io_d_out;
  wire  _T_12_io_v;
  wire  _T_13_clock;
  wire  _T_13_reset;
  wire [15:0] _T_13_io_d_in;
  wire  _T_13_io_rdy;
  wire [15:0] _T_13_io_d_out;
  wire  _T_13_io_v;
  wire  _T_14_clock;
  wire  _T_14_reset;
  wire [15:0] _T_14_io_d_in;
  wire  _T_14_io_rdy;
  wire [15:0] _T_14_io_d_out;
  wire  _T_14_io_v;
  wire  _T_15_clock;
  wire  _T_15_reset;
  wire [15:0] _T_15_io_d_in;
  wire  _T_15_io_rdy;
  wire [15:0] _T_15_io_d_out;
  wire  _T_15_io_v;
  wire  _T_16;
  wire  _T_17;
  wire  _T_18;
  wire  _T_19;
  wire  _T_20;
  wire  _T_21;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_26;
  wire  _T_27;
  wire  _T_28;
  wire  _T_29;
  MaxPool1 _T (
    .clock(_T_clock),
    .reset(_T_reset),
    .io_d_in(_T_io_d_in),
    .io_rdy(_T_io_rdy),
    .io_d_out(_T_io_d_out),
    .io_v(_T_io_v)
  );
  MaxPool1 _T_1 (
    .clock(_T_1_clock),
    .reset(_T_1_reset),
    .io_d_in(_T_1_io_d_in),
    .io_rdy(_T_1_io_rdy),
    .io_d_out(_T_1_io_d_out),
    .io_v(_T_1_io_v)
  );
  MaxPool1 _T_2 (
    .clock(_T_2_clock),
    .reset(_T_2_reset),
    .io_d_in(_T_2_io_d_in),
    .io_rdy(_T_2_io_rdy),
    .io_d_out(_T_2_io_d_out),
    .io_v(_T_2_io_v)
  );
  MaxPool1 _T_3 (
    .clock(_T_3_clock),
    .reset(_T_3_reset),
    .io_d_in(_T_3_io_d_in),
    .io_rdy(_T_3_io_rdy),
    .io_d_out(_T_3_io_d_out),
    .io_v(_T_3_io_v)
  );
  MaxPool1 _T_4 (
    .clock(_T_4_clock),
    .reset(_T_4_reset),
    .io_d_in(_T_4_io_d_in),
    .io_rdy(_T_4_io_rdy),
    .io_d_out(_T_4_io_d_out),
    .io_v(_T_4_io_v)
  );
  MaxPool1 _T_5 (
    .clock(_T_5_clock),
    .reset(_T_5_reset),
    .io_d_in(_T_5_io_d_in),
    .io_rdy(_T_5_io_rdy),
    .io_d_out(_T_5_io_d_out),
    .io_v(_T_5_io_v)
  );
  MaxPool1 _T_6 (
    .clock(_T_6_clock),
    .reset(_T_6_reset),
    .io_d_in(_T_6_io_d_in),
    .io_rdy(_T_6_io_rdy),
    .io_d_out(_T_6_io_d_out),
    .io_v(_T_6_io_v)
  );
  MaxPool1 _T_7 (
    .clock(_T_7_clock),
    .reset(_T_7_reset),
    .io_d_in(_T_7_io_d_in),
    .io_rdy(_T_7_io_rdy),
    .io_d_out(_T_7_io_d_out),
    .io_v(_T_7_io_v)
  );
  MaxPool1 _T_8 (
    .clock(_T_8_clock),
    .reset(_T_8_reset),
    .io_d_in(_T_8_io_d_in),
    .io_rdy(_T_8_io_rdy),
    .io_d_out(_T_8_io_d_out),
    .io_v(_T_8_io_v)
  );
  MaxPool1 _T_9 (
    .clock(_T_9_clock),
    .reset(_T_9_reset),
    .io_d_in(_T_9_io_d_in),
    .io_rdy(_T_9_io_rdy),
    .io_d_out(_T_9_io_d_out),
    .io_v(_T_9_io_v)
  );
  MaxPool1 _T_10 (
    .clock(_T_10_clock),
    .reset(_T_10_reset),
    .io_d_in(_T_10_io_d_in),
    .io_rdy(_T_10_io_rdy),
    .io_d_out(_T_10_io_d_out),
    .io_v(_T_10_io_v)
  );
  MaxPool1 _T_11 (
    .clock(_T_11_clock),
    .reset(_T_11_reset),
    .io_d_in(_T_11_io_d_in),
    .io_rdy(_T_11_io_rdy),
    .io_d_out(_T_11_io_d_out),
    .io_v(_T_11_io_v)
  );
  MaxPool1 _T_12 (
    .clock(_T_12_clock),
    .reset(_T_12_reset),
    .io_d_in(_T_12_io_d_in),
    .io_rdy(_T_12_io_rdy),
    .io_d_out(_T_12_io_d_out),
    .io_v(_T_12_io_v)
  );
  MaxPool1 _T_13 (
    .clock(_T_13_clock),
    .reset(_T_13_reset),
    .io_d_in(_T_13_io_d_in),
    .io_rdy(_T_13_io_rdy),
    .io_d_out(_T_13_io_d_out),
    .io_v(_T_13_io_v)
  );
  MaxPool1 _T_14 (
    .clock(_T_14_clock),
    .reset(_T_14_reset),
    .io_d_in(_T_14_io_d_in),
    .io_rdy(_T_14_io_rdy),
    .io_d_out(_T_14_io_d_out),
    .io_v(_T_14_io_v)
  );
  MaxPool1 _T_15 (
    .clock(_T_15_clock),
    .reset(_T_15_reset),
    .io_d_in(_T_15_io_d_in),
    .io_rdy(_T_15_io_rdy),
    .io_d_out(_T_15_io_d_out),
    .io_v(_T_15_io_v)
  );
  assign _T_16 = _T_io_v & _T_1_io_v;
  assign _T_17 = _T_16 & _T_2_io_v;
  assign _T_18 = _T_17 & _T_3_io_v;
  assign _T_19 = _T_18 & _T_4_io_v;
  assign _T_20 = _T_19 & _T_5_io_v;
  assign _T_21 = _T_20 & _T_6_io_v;
  assign _T_22 = _T_21 & _T_7_io_v;
  assign _T_23 = _T_22 & _T_8_io_v;
  assign _T_24 = _T_23 & _T_9_io_v;
  assign _T_25 = _T_24 & _T_10_io_v;
  assign _T_26 = _T_25 & _T_11_io_v;
  assign _T_27 = _T_26 & _T_12_io_v;
  assign _T_28 = _T_27 & _T_13_io_v;
  assign _T_29 = _T_28 & _T_14_io_v;
  assign io_d_out_0 = _T_io_d_out;
  assign io_d_out_1 = _T_1_io_d_out;
  assign io_d_out_2 = _T_2_io_d_out;
  assign io_d_out_3 = _T_3_io_d_out;
  assign io_d_out_4 = _T_4_io_d_out;
  assign io_d_out_5 = _T_5_io_d_out;
  assign io_d_out_6 = _T_6_io_d_out;
  assign io_d_out_7 = _T_7_io_d_out;
  assign io_d_out_8 = _T_8_io_d_out;
  assign io_d_out_9 = _T_9_io_d_out;
  assign io_d_out_10 = _T_10_io_d_out;
  assign io_d_out_11 = _T_11_io_d_out;
  assign io_d_out_12 = _T_12_io_d_out;
  assign io_d_out_13 = _T_13_io_d_out;
  assign io_d_out_14 = _T_14_io_d_out;
  assign io_d_out_15 = _T_15_io_d_out;
  assign io_pool_v = _T_29 & _T_15_io_v;
  assign _T_clock = clock;
  assign _T_reset = reset;
  assign _T_io_d_in = io_d_in_0;
  assign _T_io_rdy = io_rdy;
  assign _T_1_clock = clock;
  assign _T_1_reset = reset;
  assign _T_1_io_d_in = io_d_in_1;
  assign _T_1_io_rdy = io_rdy;
  assign _T_2_clock = clock;
  assign _T_2_reset = reset;
  assign _T_2_io_d_in = io_d_in_2;
  assign _T_2_io_rdy = io_rdy;
  assign _T_3_clock = clock;
  assign _T_3_reset = reset;
  assign _T_3_io_d_in = io_d_in_3;
  assign _T_3_io_rdy = io_rdy;
  assign _T_4_clock = clock;
  assign _T_4_reset = reset;
  assign _T_4_io_d_in = io_d_in_4;
  assign _T_4_io_rdy = io_rdy;
  assign _T_5_clock = clock;
  assign _T_5_reset = reset;
  assign _T_5_io_d_in = io_d_in_5;
  assign _T_5_io_rdy = io_rdy;
  assign _T_6_clock = clock;
  assign _T_6_reset = reset;
  assign _T_6_io_d_in = io_d_in_6;
  assign _T_6_io_rdy = io_rdy;
  assign _T_7_clock = clock;
  assign _T_7_reset = reset;
  assign _T_7_io_d_in = io_d_in_7;
  assign _T_7_io_rdy = io_rdy;
  assign _T_8_clock = clock;
  assign _T_8_reset = reset;
  assign _T_8_io_d_in = io_d_in_8;
  assign _T_8_io_rdy = io_rdy;
  assign _T_9_clock = clock;
  assign _T_9_reset = reset;
  assign _T_9_io_d_in = io_d_in_9;
  assign _T_9_io_rdy = io_rdy;
  assign _T_10_clock = clock;
  assign _T_10_reset = reset;
  assign _T_10_io_d_in = io_d_in_10;
  assign _T_10_io_rdy = io_rdy;
  assign _T_11_clock = clock;
  assign _T_11_reset = reset;
  assign _T_11_io_d_in = io_d_in_11;
  assign _T_11_io_rdy = io_rdy;
  assign _T_12_clock = clock;
  assign _T_12_reset = reset;
  assign _T_12_io_d_in = io_d_in_12;
  assign _T_12_io_rdy = io_rdy;
  assign _T_13_clock = clock;
  assign _T_13_reset = reset;
  assign _T_13_io_d_in = io_d_in_13;
  assign _T_13_io_rdy = io_rdy;
  assign _T_14_clock = clock;
  assign _T_14_reset = reset;
  assign _T_14_io_d_in = io_d_in_14;
  assign _T_14_io_rdy = io_rdy;
  assign _T_15_clock = clock;
  assign _T_15_reset = reset;
  assign _T_15_io_d_in = io_d_in_15;
  assign _T_15_io_rdy = io_rdy;
endmodule
module Mac_102(
  input           clock,
  input           reset,
  input  [6399:0] io_a,
  input  [6399:0] io_b,
  input           io_rdy,
  output [31:0]   io_q,
  output          io_v
);
  wire [15:0] a_0;
  wire [15:0] b_0;
  wire [15:0] a_1;
  wire [15:0] b_1;
  wire [15:0] a_2;
  wire [15:0] b_2;
  wire [15:0] a_3;
  wire [15:0] b_3;
  wire [15:0] a_4;
  wire [15:0] b_4;
  wire [15:0] a_5;
  wire [15:0] b_5;
  wire [15:0] a_6;
  wire [15:0] b_6;
  wire [15:0] a_7;
  wire [15:0] b_7;
  wire [15:0] a_8;
  wire [15:0] b_8;
  wire [15:0] a_9;
  wire [15:0] b_9;
  wire [15:0] a_10;
  wire [15:0] b_10;
  wire [15:0] a_11;
  wire [15:0] b_11;
  wire [15:0] a_12;
  wire [15:0] b_12;
  wire [15:0] a_13;
  wire [15:0] b_13;
  wire [15:0] a_14;
  wire [15:0] b_14;
  wire [15:0] a_15;
  wire [15:0] b_15;
  wire [15:0] a_16;
  wire [15:0] b_16;
  wire [15:0] a_17;
  wire [15:0] b_17;
  wire [15:0] a_18;
  wire [15:0] b_18;
  wire [15:0] a_19;
  wire [15:0] b_19;
  wire [15:0] a_20;
  wire [15:0] b_20;
  wire [15:0] a_21;
  wire [15:0] b_21;
  wire [15:0] a_22;
  wire [15:0] b_22;
  wire [15:0] a_23;
  wire [15:0] b_23;
  wire [15:0] a_24;
  wire [15:0] b_24;
  wire [15:0] a_25;
  wire [15:0] b_25;
  wire [15:0] a_26;
  wire [15:0] b_26;
  wire [15:0] a_27;
  wire [15:0] b_27;
  wire [15:0] a_28;
  wire [15:0] b_28;
  wire [15:0] a_29;
  wire [15:0] b_29;
  wire [15:0] a_30;
  wire [15:0] b_30;
  wire [15:0] a_31;
  wire [15:0] b_31;
  wire [15:0] a_32;
  wire [15:0] b_32;
  wire [15:0] a_33;
  wire [15:0] b_33;
  wire [15:0] a_34;
  wire [15:0] b_34;
  wire [15:0] a_35;
  wire [15:0] b_35;
  wire [15:0] a_36;
  wire [15:0] b_36;
  wire [15:0] a_37;
  wire [15:0] b_37;
  wire [15:0] a_38;
  wire [15:0] b_38;
  wire [15:0] a_39;
  wire [15:0] b_39;
  wire [15:0] a_40;
  wire [15:0] b_40;
  wire [15:0] a_41;
  wire [15:0] b_41;
  wire [15:0] a_42;
  wire [15:0] b_42;
  wire [15:0] a_43;
  wire [15:0] b_43;
  wire [15:0] a_44;
  wire [15:0] b_44;
  wire [15:0] a_45;
  wire [15:0] b_45;
  wire [15:0] a_46;
  wire [15:0] b_46;
  wire [15:0] a_47;
  wire [15:0] b_47;
  wire [15:0] a_48;
  wire [15:0] b_48;
  wire [15:0] a_49;
  wire [15:0] b_49;
  wire [15:0] a_50;
  wire [15:0] b_50;
  wire [15:0] a_51;
  wire [15:0] b_51;
  wire [15:0] a_52;
  wire [15:0] b_52;
  wire [15:0] a_53;
  wire [15:0] b_53;
  wire [15:0] a_54;
  wire [15:0] b_54;
  wire [15:0] a_55;
  wire [15:0] b_55;
  wire [15:0] a_56;
  wire [15:0] b_56;
  wire [15:0] a_57;
  wire [15:0] b_57;
  wire [15:0] a_58;
  wire [15:0] b_58;
  wire [15:0] a_59;
  wire [15:0] b_59;
  wire [15:0] a_60;
  wire [15:0] b_60;
  wire [15:0] a_61;
  wire [15:0] b_61;
  wire [15:0] a_62;
  wire [15:0] b_62;
  wire [15:0] a_63;
  wire [15:0] b_63;
  wire [15:0] a_64;
  wire [15:0] b_64;
  wire [15:0] a_65;
  wire [15:0] b_65;
  wire [15:0] a_66;
  wire [15:0] b_66;
  wire [15:0] a_67;
  wire [15:0] b_67;
  wire [15:0] a_68;
  wire [15:0] b_68;
  wire [15:0] a_69;
  wire [15:0] b_69;
  wire [15:0] a_70;
  wire [15:0] b_70;
  wire [15:0] a_71;
  wire [15:0] b_71;
  wire [15:0] a_72;
  wire [15:0] b_72;
  wire [15:0] a_73;
  wire [15:0] b_73;
  wire [15:0] a_74;
  wire [15:0] b_74;
  wire [15:0] a_75;
  wire [15:0] b_75;
  wire [15:0] a_76;
  wire [15:0] b_76;
  wire [15:0] a_77;
  wire [15:0] b_77;
  wire [15:0] a_78;
  wire [15:0] b_78;
  wire [15:0] a_79;
  wire [15:0] b_79;
  wire [15:0] a_80;
  wire [15:0] b_80;
  wire [15:0] a_81;
  wire [15:0] b_81;
  wire [15:0] a_82;
  wire [15:0] b_82;
  wire [15:0] a_83;
  wire [15:0] b_83;
  wire [15:0] a_84;
  wire [15:0] b_84;
  wire [15:0] a_85;
  wire [15:0] b_85;
  wire [15:0] a_86;
  wire [15:0] b_86;
  wire [15:0] a_87;
  wire [15:0] b_87;
  wire [15:0] a_88;
  wire [15:0] b_88;
  wire [15:0] a_89;
  wire [15:0] b_89;
  wire [15:0] a_90;
  wire [15:0] b_90;
  wire [15:0] a_91;
  wire [15:0] b_91;
  wire [15:0] a_92;
  wire [15:0] b_92;
  wire [15:0] a_93;
  wire [15:0] b_93;
  wire [15:0] a_94;
  wire [15:0] b_94;
  wire [15:0] a_95;
  wire [15:0] b_95;
  wire [15:0] a_96;
  wire [15:0] b_96;
  wire [15:0] a_97;
  wire [15:0] b_97;
  wire [15:0] a_98;
  wire [15:0] b_98;
  wire [15:0] a_99;
  wire [15:0] b_99;
  wire [15:0] a_100;
  wire [15:0] b_100;
  wire [15:0] a_101;
  wire [15:0] b_101;
  wire [15:0] a_102;
  wire [15:0] b_102;
  wire [15:0] a_103;
  wire [15:0] b_103;
  wire [15:0] a_104;
  wire [15:0] b_104;
  wire [15:0] a_105;
  wire [15:0] b_105;
  wire [15:0] a_106;
  wire [15:0] b_106;
  wire [15:0] a_107;
  wire [15:0] b_107;
  wire [15:0] a_108;
  wire [15:0] b_108;
  wire [15:0] a_109;
  wire [15:0] b_109;
  wire [15:0] a_110;
  wire [15:0] b_110;
  wire [15:0] a_111;
  wire [15:0] b_111;
  wire [15:0] a_112;
  wire [15:0] b_112;
  wire [15:0] a_113;
  wire [15:0] b_113;
  wire [15:0] a_114;
  wire [15:0] b_114;
  wire [15:0] a_115;
  wire [15:0] b_115;
  wire [15:0] a_116;
  wire [15:0] b_116;
  wire [15:0] a_117;
  wire [15:0] b_117;
  wire [15:0] a_118;
  wire [15:0] b_118;
  wire [15:0] a_119;
  wire [15:0] b_119;
  wire [15:0] a_120;
  wire [15:0] b_120;
  wire [15:0] a_121;
  wire [15:0] b_121;
  wire [15:0] a_122;
  wire [15:0] b_122;
  wire [15:0] a_123;
  wire [15:0] b_123;
  wire [15:0] a_124;
  wire [15:0] b_124;
  wire [15:0] a_125;
  wire [15:0] b_125;
  wire [15:0] a_126;
  wire [15:0] b_126;
  wire [15:0] a_127;
  wire [15:0] b_127;
  wire [15:0] a_128;
  wire [15:0] b_128;
  wire [15:0] a_129;
  wire [15:0] b_129;
  wire [15:0] a_130;
  wire [15:0] b_130;
  wire [15:0] a_131;
  wire [15:0] b_131;
  wire [15:0] a_132;
  wire [15:0] b_132;
  wire [15:0] a_133;
  wire [15:0] b_133;
  wire [15:0] a_134;
  wire [15:0] b_134;
  wire [15:0] a_135;
  wire [15:0] b_135;
  wire [15:0] a_136;
  wire [15:0] b_136;
  wire [15:0] a_137;
  wire [15:0] b_137;
  wire [15:0] a_138;
  wire [15:0] b_138;
  wire [15:0] a_139;
  wire [15:0] b_139;
  wire [15:0] a_140;
  wire [15:0] b_140;
  wire [15:0] a_141;
  wire [15:0] b_141;
  wire [15:0] a_142;
  wire [15:0] b_142;
  wire [15:0] a_143;
  wire [15:0] b_143;
  wire [15:0] a_144;
  wire [15:0] b_144;
  wire [15:0] a_145;
  wire [15:0] b_145;
  wire [15:0] a_146;
  wire [15:0] b_146;
  wire [15:0] a_147;
  wire [15:0] b_147;
  wire [15:0] a_148;
  wire [15:0] b_148;
  wire [15:0] a_149;
  wire [15:0] b_149;
  wire [15:0] a_150;
  wire [15:0] b_150;
  wire [15:0] a_151;
  wire [15:0] b_151;
  wire [15:0] a_152;
  wire [15:0] b_152;
  wire [15:0] a_153;
  wire [15:0] b_153;
  wire [15:0] a_154;
  wire [15:0] b_154;
  wire [15:0] a_155;
  wire [15:0] b_155;
  wire [15:0] a_156;
  wire [15:0] b_156;
  wire [15:0] a_157;
  wire [15:0] b_157;
  wire [15:0] a_158;
  wire [15:0] b_158;
  wire [15:0] a_159;
  wire [15:0] b_159;
  wire [15:0] a_160;
  wire [15:0] b_160;
  wire [15:0] a_161;
  wire [15:0] b_161;
  wire [15:0] a_162;
  wire [15:0] b_162;
  wire [15:0] a_163;
  wire [15:0] b_163;
  wire [15:0] a_164;
  wire [15:0] b_164;
  wire [15:0] a_165;
  wire [15:0] b_165;
  wire [15:0] a_166;
  wire [15:0] b_166;
  wire [15:0] a_167;
  wire [15:0] b_167;
  wire [15:0] a_168;
  wire [15:0] b_168;
  wire [15:0] a_169;
  wire [15:0] b_169;
  wire [15:0] a_170;
  wire [15:0] b_170;
  wire [15:0] a_171;
  wire [15:0] b_171;
  wire [15:0] a_172;
  wire [15:0] b_172;
  wire [15:0] a_173;
  wire [15:0] b_173;
  wire [15:0] a_174;
  wire [15:0] b_174;
  wire [15:0] a_175;
  wire [15:0] b_175;
  wire [15:0] a_176;
  wire [15:0] b_176;
  wire [15:0] a_177;
  wire [15:0] b_177;
  wire [15:0] a_178;
  wire [15:0] b_178;
  wire [15:0] a_179;
  wire [15:0] b_179;
  wire [15:0] a_180;
  wire [15:0] b_180;
  wire [15:0] a_181;
  wire [15:0] b_181;
  wire [15:0] a_182;
  wire [15:0] b_182;
  wire [15:0] a_183;
  wire [15:0] b_183;
  wire [15:0] a_184;
  wire [15:0] b_184;
  wire [15:0] a_185;
  wire [15:0] b_185;
  wire [15:0] a_186;
  wire [15:0] b_186;
  wire [15:0] a_187;
  wire [15:0] b_187;
  wire [15:0] a_188;
  wire [15:0] b_188;
  wire [15:0] a_189;
  wire [15:0] b_189;
  wire [15:0] a_190;
  wire [15:0] b_190;
  wire [15:0] a_191;
  wire [15:0] b_191;
  wire [15:0] a_192;
  wire [15:0] b_192;
  wire [15:0] a_193;
  wire [15:0] b_193;
  wire [15:0] a_194;
  wire [15:0] b_194;
  wire [15:0] a_195;
  wire [15:0] b_195;
  wire [15:0] a_196;
  wire [15:0] b_196;
  wire [15:0] a_197;
  wire [15:0] b_197;
  wire [15:0] a_198;
  wire [15:0] b_198;
  wire [15:0] a_199;
  wire [15:0] b_199;
  wire [15:0] a_200;
  wire [15:0] b_200;
  wire [15:0] a_201;
  wire [15:0] b_201;
  wire [15:0] a_202;
  wire [15:0] b_202;
  wire [15:0] a_203;
  wire [15:0] b_203;
  wire [15:0] a_204;
  wire [15:0] b_204;
  wire [15:0] a_205;
  wire [15:0] b_205;
  wire [15:0] a_206;
  wire [15:0] b_206;
  wire [15:0] a_207;
  wire [15:0] b_207;
  wire [15:0] a_208;
  wire [15:0] b_208;
  wire [15:0] a_209;
  wire [15:0] b_209;
  wire [15:0] a_210;
  wire [15:0] b_210;
  wire [15:0] a_211;
  wire [15:0] b_211;
  wire [15:0] a_212;
  wire [15:0] b_212;
  wire [15:0] a_213;
  wire [15:0] b_213;
  wire [15:0] a_214;
  wire [15:0] b_214;
  wire [15:0] a_215;
  wire [15:0] b_215;
  wire [15:0] a_216;
  wire [15:0] b_216;
  wire [15:0] a_217;
  wire [15:0] b_217;
  wire [15:0] a_218;
  wire [15:0] b_218;
  wire [15:0] a_219;
  wire [15:0] b_219;
  wire [15:0] a_220;
  wire [15:0] b_220;
  wire [15:0] a_221;
  wire [15:0] b_221;
  wire [15:0] a_222;
  wire [15:0] b_222;
  wire [15:0] a_223;
  wire [15:0] b_223;
  wire [15:0] a_224;
  wire [15:0] b_224;
  wire [15:0] a_225;
  wire [15:0] b_225;
  wire [15:0] a_226;
  wire [15:0] b_226;
  wire [15:0] a_227;
  wire [15:0] b_227;
  wire [15:0] a_228;
  wire [15:0] b_228;
  wire [15:0] a_229;
  wire [15:0] b_229;
  wire [15:0] a_230;
  wire [15:0] b_230;
  wire [15:0] a_231;
  wire [15:0] b_231;
  wire [15:0] a_232;
  wire [15:0] b_232;
  wire [15:0] a_233;
  wire [15:0] b_233;
  wire [15:0] a_234;
  wire [15:0] b_234;
  wire [15:0] a_235;
  wire [15:0] b_235;
  wire [15:0] a_236;
  wire [15:0] b_236;
  wire [15:0] a_237;
  wire [15:0] b_237;
  wire [15:0] a_238;
  wire [15:0] b_238;
  wire [15:0] a_239;
  wire [15:0] b_239;
  wire [15:0] a_240;
  wire [15:0] b_240;
  wire [15:0] a_241;
  wire [15:0] b_241;
  wire [15:0] a_242;
  wire [15:0] b_242;
  wire [15:0] a_243;
  wire [15:0] b_243;
  wire [15:0] a_244;
  wire [15:0] b_244;
  wire [15:0] a_245;
  wire [15:0] b_245;
  wire [15:0] a_246;
  wire [15:0] b_246;
  wire [15:0] a_247;
  wire [15:0] b_247;
  wire [15:0] a_248;
  wire [15:0] b_248;
  wire [15:0] a_249;
  wire [15:0] b_249;
  wire [15:0] a_250;
  wire [15:0] b_250;
  wire [15:0] a_251;
  wire [15:0] b_251;
  wire [15:0] a_252;
  wire [15:0] b_252;
  wire [15:0] a_253;
  wire [15:0] b_253;
  wire [15:0] a_254;
  wire [15:0] b_254;
  wire [15:0] a_255;
  wire [15:0] b_255;
  wire [15:0] a_256;
  wire [15:0] b_256;
  wire [15:0] a_257;
  wire [15:0] b_257;
  wire [15:0] a_258;
  wire [15:0] b_258;
  wire [15:0] a_259;
  wire [15:0] b_259;
  wire [15:0] a_260;
  wire [15:0] b_260;
  wire [15:0] a_261;
  wire [15:0] b_261;
  wire [15:0] a_262;
  wire [15:0] b_262;
  wire [15:0] a_263;
  wire [15:0] b_263;
  wire [15:0] a_264;
  wire [15:0] b_264;
  wire [15:0] a_265;
  wire [15:0] b_265;
  wire [15:0] a_266;
  wire [15:0] b_266;
  wire [15:0] a_267;
  wire [15:0] b_267;
  wire [15:0] a_268;
  wire [15:0] b_268;
  wire [15:0] a_269;
  wire [15:0] b_269;
  wire [15:0] a_270;
  wire [15:0] b_270;
  wire [15:0] a_271;
  wire [15:0] b_271;
  wire [15:0] a_272;
  wire [15:0] b_272;
  wire [15:0] a_273;
  wire [15:0] b_273;
  wire [15:0] a_274;
  wire [15:0] b_274;
  wire [15:0] a_275;
  wire [15:0] b_275;
  wire [15:0] a_276;
  wire [15:0] b_276;
  wire [15:0] a_277;
  wire [15:0] b_277;
  wire [15:0] a_278;
  wire [15:0] b_278;
  wire [15:0] a_279;
  wire [15:0] b_279;
  wire [15:0] a_280;
  wire [15:0] b_280;
  wire [15:0] a_281;
  wire [15:0] b_281;
  wire [15:0] a_282;
  wire [15:0] b_282;
  wire [15:0] a_283;
  wire [15:0] b_283;
  wire [15:0] a_284;
  wire [15:0] b_284;
  wire [15:0] a_285;
  wire [15:0] b_285;
  wire [15:0] a_286;
  wire [15:0] b_286;
  wire [15:0] a_287;
  wire [15:0] b_287;
  wire [15:0] a_288;
  wire [15:0] b_288;
  wire [15:0] a_289;
  wire [15:0] b_289;
  wire [15:0] a_290;
  wire [15:0] b_290;
  wire [15:0] a_291;
  wire [15:0] b_291;
  wire [15:0] a_292;
  wire [15:0] b_292;
  wire [15:0] a_293;
  wire [15:0] b_293;
  wire [15:0] a_294;
  wire [15:0] b_294;
  wire [15:0] a_295;
  wire [15:0] b_295;
  wire [15:0] a_296;
  wire [15:0] b_296;
  wire [15:0] a_297;
  wire [15:0] b_297;
  wire [15:0] a_298;
  wire [15:0] b_298;
  wire [15:0] a_299;
  wire [15:0] b_299;
  wire [15:0] a_300;
  wire [15:0] b_300;
  wire [15:0] a_301;
  wire [15:0] b_301;
  wire [15:0] a_302;
  wire [15:0] b_302;
  wire [15:0] a_303;
  wire [15:0] b_303;
  wire [15:0] a_304;
  wire [15:0] b_304;
  wire [15:0] a_305;
  wire [15:0] b_305;
  wire [15:0] a_306;
  wire [15:0] b_306;
  wire [15:0] a_307;
  wire [15:0] b_307;
  wire [15:0] a_308;
  wire [15:0] b_308;
  wire [15:0] a_309;
  wire [15:0] b_309;
  wire [15:0] a_310;
  wire [15:0] b_310;
  wire [15:0] a_311;
  wire [15:0] b_311;
  wire [15:0] a_312;
  wire [15:0] b_312;
  wire [15:0] a_313;
  wire [15:0] b_313;
  wire [15:0] a_314;
  wire [15:0] b_314;
  wire [15:0] a_315;
  wire [15:0] b_315;
  wire [15:0] a_316;
  wire [15:0] b_316;
  wire [15:0] a_317;
  wire [15:0] b_317;
  wire [15:0] a_318;
  wire [15:0] b_318;
  wire [15:0] a_319;
  wire [15:0] b_319;
  wire [15:0] a_320;
  wire [15:0] b_320;
  wire [15:0] a_321;
  wire [15:0] b_321;
  wire [15:0] a_322;
  wire [15:0] b_322;
  wire [15:0] a_323;
  wire [15:0] b_323;
  wire [15:0] a_324;
  wire [15:0] b_324;
  wire [15:0] a_325;
  wire [15:0] b_325;
  wire [15:0] a_326;
  wire [15:0] b_326;
  wire [15:0] a_327;
  wire [15:0] b_327;
  wire [15:0] a_328;
  wire [15:0] b_328;
  wire [15:0] a_329;
  wire [15:0] b_329;
  wire [15:0] a_330;
  wire [15:0] b_330;
  wire [15:0] a_331;
  wire [15:0] b_331;
  wire [15:0] a_332;
  wire [15:0] b_332;
  wire [15:0] a_333;
  wire [15:0] b_333;
  wire [15:0] a_334;
  wire [15:0] b_334;
  wire [15:0] a_335;
  wire [15:0] b_335;
  wire [15:0] a_336;
  wire [15:0] b_336;
  wire [15:0] a_337;
  wire [15:0] b_337;
  wire [15:0] a_338;
  wire [15:0] b_338;
  wire [15:0] a_339;
  wire [15:0] b_339;
  wire [15:0] a_340;
  wire [15:0] b_340;
  wire [15:0] a_341;
  wire [15:0] b_341;
  wire [15:0] a_342;
  wire [15:0] b_342;
  wire [15:0] a_343;
  wire [15:0] b_343;
  wire [15:0] a_344;
  wire [15:0] b_344;
  wire [15:0] a_345;
  wire [15:0] b_345;
  wire [15:0] a_346;
  wire [15:0] b_346;
  wire [15:0] a_347;
  wire [15:0] b_347;
  wire [15:0] a_348;
  wire [15:0] b_348;
  wire [15:0] a_349;
  wire [15:0] b_349;
  wire [15:0] a_350;
  wire [15:0] b_350;
  wire [15:0] a_351;
  wire [15:0] b_351;
  wire [15:0] a_352;
  wire [15:0] b_352;
  wire [15:0] a_353;
  wire [15:0] b_353;
  wire [15:0] a_354;
  wire [15:0] b_354;
  wire [15:0] a_355;
  wire [15:0] b_355;
  wire [15:0] a_356;
  wire [15:0] b_356;
  wire [15:0] a_357;
  wire [15:0] b_357;
  wire [15:0] a_358;
  wire [15:0] b_358;
  wire [15:0] a_359;
  wire [15:0] b_359;
  wire [15:0] a_360;
  wire [15:0] b_360;
  wire [15:0] a_361;
  wire [15:0] b_361;
  wire [15:0] a_362;
  wire [15:0] b_362;
  wire [15:0] a_363;
  wire [15:0] b_363;
  wire [15:0] a_364;
  wire [15:0] b_364;
  wire [15:0] a_365;
  wire [15:0] b_365;
  wire [15:0] a_366;
  wire [15:0] b_366;
  wire [15:0] a_367;
  wire [15:0] b_367;
  wire [15:0] a_368;
  wire [15:0] b_368;
  wire [15:0] a_369;
  wire [15:0] b_369;
  wire [15:0] a_370;
  wire [15:0] b_370;
  wire [15:0] a_371;
  wire [15:0] b_371;
  wire [15:0] a_372;
  wire [15:0] b_372;
  wire [15:0] a_373;
  wire [15:0] b_373;
  wire [15:0] a_374;
  wire [15:0] b_374;
  wire [15:0] a_375;
  wire [15:0] b_375;
  wire [15:0] a_376;
  wire [15:0] b_376;
  wire [15:0] a_377;
  wire [15:0] b_377;
  wire [15:0] a_378;
  wire [15:0] b_378;
  wire [15:0] a_379;
  wire [15:0] b_379;
  wire [15:0] a_380;
  wire [15:0] b_380;
  wire [15:0] a_381;
  wire [15:0] b_381;
  wire [15:0] a_382;
  wire [15:0] b_382;
  wire [15:0] a_383;
  wire [15:0] b_383;
  wire [15:0] a_384;
  wire [15:0] b_384;
  wire [15:0] a_385;
  wire [15:0] b_385;
  wire [15:0] a_386;
  wire [15:0] b_386;
  wire [15:0] a_387;
  wire [15:0] b_387;
  wire [15:0] a_388;
  wire [15:0] b_388;
  wire [15:0] a_389;
  wire [15:0] b_389;
  wire [15:0] a_390;
  wire [15:0] b_390;
  wire [15:0] a_391;
  wire [15:0] b_391;
  wire [15:0] a_392;
  wire [15:0] b_392;
  wire [15:0] a_393;
  wire [15:0] b_393;
  wire [15:0] a_394;
  wire [15:0] b_394;
  wire [15:0] a_395;
  wire [15:0] b_395;
  wire [15:0] a_396;
  wire [15:0] b_396;
  wire [15:0] a_397;
  wire [15:0] b_397;
  wire [15:0] a_398;
  wire [15:0] b_398;
  wire [15:0] a_399;
  wire [15:0] b_399;
  reg [31:0] sum;
  reg [31:0] _RAND_0;
  reg [8:0] i;
  reg [31:0] _RAND_1;
  wire  _T_803;
  wire  _T_804;
  wire [15:0] _GEN_1;
  wire [15:0] _GEN_2;
  wire [15:0] _GEN_3;
  wire [15:0] _GEN_4;
  wire [15:0] _GEN_5;
  wire [15:0] _GEN_6;
  wire [15:0] _GEN_7;
  wire [15:0] _GEN_8;
  wire [15:0] _GEN_9;
  wire [15:0] _GEN_10;
  wire [15:0] _GEN_11;
  wire [15:0] _GEN_12;
  wire [15:0] _GEN_13;
  wire [15:0] _GEN_14;
  wire [15:0] _GEN_15;
  wire [15:0] _GEN_16;
  wire [15:0] _GEN_17;
  wire [15:0] _GEN_18;
  wire [15:0] _GEN_19;
  wire [15:0] _GEN_20;
  wire [15:0] _GEN_21;
  wire [15:0] _GEN_22;
  wire [15:0] _GEN_23;
  wire [15:0] _GEN_24;
  wire [15:0] _GEN_25;
  wire [15:0] _GEN_26;
  wire [15:0] _GEN_27;
  wire [15:0] _GEN_28;
  wire [15:0] _GEN_29;
  wire [15:0] _GEN_30;
  wire [15:0] _GEN_31;
  wire [15:0] _GEN_32;
  wire [15:0] _GEN_33;
  wire [15:0] _GEN_34;
  wire [15:0] _GEN_35;
  wire [15:0] _GEN_36;
  wire [15:0] _GEN_37;
  wire [15:0] _GEN_38;
  wire [15:0] _GEN_39;
  wire [15:0] _GEN_40;
  wire [15:0] _GEN_41;
  wire [15:0] _GEN_42;
  wire [15:0] _GEN_43;
  wire [15:0] _GEN_44;
  wire [15:0] _GEN_45;
  wire [15:0] _GEN_46;
  wire [15:0] _GEN_47;
  wire [15:0] _GEN_48;
  wire [15:0] _GEN_49;
  wire [15:0] _GEN_50;
  wire [15:0] _GEN_51;
  wire [15:0] _GEN_52;
  wire [15:0] _GEN_53;
  wire [15:0] _GEN_54;
  wire [15:0] _GEN_55;
  wire [15:0] _GEN_56;
  wire [15:0] _GEN_57;
  wire [15:0] _GEN_58;
  wire [15:0] _GEN_59;
  wire [15:0] _GEN_60;
  wire [15:0] _GEN_61;
  wire [15:0] _GEN_62;
  wire [15:0] _GEN_63;
  wire [15:0] _GEN_64;
  wire [15:0] _GEN_65;
  wire [15:0] _GEN_66;
  wire [15:0] _GEN_67;
  wire [15:0] _GEN_68;
  wire [15:0] _GEN_69;
  wire [15:0] _GEN_70;
  wire [15:0] _GEN_71;
  wire [15:0] _GEN_72;
  wire [15:0] _GEN_73;
  wire [15:0] _GEN_74;
  wire [15:0] _GEN_75;
  wire [15:0] _GEN_76;
  wire [15:0] _GEN_77;
  wire [15:0] _GEN_78;
  wire [15:0] _GEN_79;
  wire [15:0] _GEN_80;
  wire [15:0] _GEN_81;
  wire [15:0] _GEN_82;
  wire [15:0] _GEN_83;
  wire [15:0] _GEN_84;
  wire [15:0] _GEN_85;
  wire [15:0] _GEN_86;
  wire [15:0] _GEN_87;
  wire [15:0] _GEN_88;
  wire [15:0] _GEN_89;
  wire [15:0] _GEN_90;
  wire [15:0] _GEN_91;
  wire [15:0] _GEN_92;
  wire [15:0] _GEN_93;
  wire [15:0] _GEN_94;
  wire [15:0] _GEN_95;
  wire [15:0] _GEN_96;
  wire [15:0] _GEN_97;
  wire [15:0] _GEN_98;
  wire [15:0] _GEN_99;
  wire [15:0] _GEN_100;
  wire [15:0] _GEN_101;
  wire [15:0] _GEN_102;
  wire [15:0] _GEN_103;
  wire [15:0] _GEN_104;
  wire [15:0] _GEN_105;
  wire [15:0] _GEN_106;
  wire [15:0] _GEN_107;
  wire [15:0] _GEN_108;
  wire [15:0] _GEN_109;
  wire [15:0] _GEN_110;
  wire [15:0] _GEN_111;
  wire [15:0] _GEN_112;
  wire [15:0] _GEN_113;
  wire [15:0] _GEN_114;
  wire [15:0] _GEN_115;
  wire [15:0] _GEN_116;
  wire [15:0] _GEN_117;
  wire [15:0] _GEN_118;
  wire [15:0] _GEN_119;
  wire [15:0] _GEN_120;
  wire [15:0] _GEN_121;
  wire [15:0] _GEN_122;
  wire [15:0] _GEN_123;
  wire [15:0] _GEN_124;
  wire [15:0] _GEN_125;
  wire [15:0] _GEN_126;
  wire [15:0] _GEN_127;
  wire [15:0] _GEN_128;
  wire [15:0] _GEN_129;
  wire [15:0] _GEN_130;
  wire [15:0] _GEN_131;
  wire [15:0] _GEN_132;
  wire [15:0] _GEN_133;
  wire [15:0] _GEN_134;
  wire [15:0] _GEN_135;
  wire [15:0] _GEN_136;
  wire [15:0] _GEN_137;
  wire [15:0] _GEN_138;
  wire [15:0] _GEN_139;
  wire [15:0] _GEN_140;
  wire [15:0] _GEN_141;
  wire [15:0] _GEN_142;
  wire [15:0] _GEN_143;
  wire [15:0] _GEN_144;
  wire [15:0] _GEN_145;
  wire [15:0] _GEN_146;
  wire [15:0] _GEN_147;
  wire [15:0] _GEN_148;
  wire [15:0] _GEN_149;
  wire [15:0] _GEN_150;
  wire [15:0] _GEN_151;
  wire [15:0] _GEN_152;
  wire [15:0] _GEN_153;
  wire [15:0] _GEN_154;
  wire [15:0] _GEN_155;
  wire [15:0] _GEN_156;
  wire [15:0] _GEN_157;
  wire [15:0] _GEN_158;
  wire [15:0] _GEN_159;
  wire [15:0] _GEN_160;
  wire [15:0] _GEN_161;
  wire [15:0] _GEN_162;
  wire [15:0] _GEN_163;
  wire [15:0] _GEN_164;
  wire [15:0] _GEN_165;
  wire [15:0] _GEN_166;
  wire [15:0] _GEN_167;
  wire [15:0] _GEN_168;
  wire [15:0] _GEN_169;
  wire [15:0] _GEN_170;
  wire [15:0] _GEN_171;
  wire [15:0] _GEN_172;
  wire [15:0] _GEN_173;
  wire [15:0] _GEN_174;
  wire [15:0] _GEN_175;
  wire [15:0] _GEN_176;
  wire [15:0] _GEN_177;
  wire [15:0] _GEN_178;
  wire [15:0] _GEN_179;
  wire [15:0] _GEN_180;
  wire [15:0] _GEN_181;
  wire [15:0] _GEN_182;
  wire [15:0] _GEN_183;
  wire [15:0] _GEN_184;
  wire [15:0] _GEN_185;
  wire [15:0] _GEN_186;
  wire [15:0] _GEN_187;
  wire [15:0] _GEN_188;
  wire [15:0] _GEN_189;
  wire [15:0] _GEN_190;
  wire [15:0] _GEN_191;
  wire [15:0] _GEN_192;
  wire [15:0] _GEN_193;
  wire [15:0] _GEN_194;
  wire [15:0] _GEN_195;
  wire [15:0] _GEN_196;
  wire [15:0] _GEN_197;
  wire [15:0] _GEN_198;
  wire [15:0] _GEN_199;
  wire [15:0] _GEN_200;
  wire [15:0] _GEN_201;
  wire [15:0] _GEN_202;
  wire [15:0] _GEN_203;
  wire [15:0] _GEN_204;
  wire [15:0] _GEN_205;
  wire [15:0] _GEN_206;
  wire [15:0] _GEN_207;
  wire [15:0] _GEN_208;
  wire [15:0] _GEN_209;
  wire [15:0] _GEN_210;
  wire [15:0] _GEN_211;
  wire [15:0] _GEN_212;
  wire [15:0] _GEN_213;
  wire [15:0] _GEN_214;
  wire [15:0] _GEN_215;
  wire [15:0] _GEN_216;
  wire [15:0] _GEN_217;
  wire [15:0] _GEN_218;
  wire [15:0] _GEN_219;
  wire [15:0] _GEN_220;
  wire [15:0] _GEN_221;
  wire [15:0] _GEN_222;
  wire [15:0] _GEN_223;
  wire [15:0] _GEN_224;
  wire [15:0] _GEN_225;
  wire [15:0] _GEN_226;
  wire [15:0] _GEN_227;
  wire [15:0] _GEN_228;
  wire [15:0] _GEN_229;
  wire [15:0] _GEN_230;
  wire [15:0] _GEN_231;
  wire [15:0] _GEN_232;
  wire [15:0] _GEN_233;
  wire [15:0] _GEN_234;
  wire [15:0] _GEN_235;
  wire [15:0] _GEN_236;
  wire [15:0] _GEN_237;
  wire [15:0] _GEN_238;
  wire [15:0] _GEN_239;
  wire [15:0] _GEN_240;
  wire [15:0] _GEN_241;
  wire [15:0] _GEN_242;
  wire [15:0] _GEN_243;
  wire [15:0] _GEN_244;
  wire [15:0] _GEN_245;
  wire [15:0] _GEN_246;
  wire [15:0] _GEN_247;
  wire [15:0] _GEN_248;
  wire [15:0] _GEN_249;
  wire [15:0] _GEN_250;
  wire [15:0] _GEN_251;
  wire [15:0] _GEN_252;
  wire [15:0] _GEN_253;
  wire [15:0] _GEN_254;
  wire [15:0] _GEN_255;
  wire [15:0] _GEN_256;
  wire [15:0] _GEN_257;
  wire [15:0] _GEN_258;
  wire [15:0] _GEN_259;
  wire [15:0] _GEN_260;
  wire [15:0] _GEN_261;
  wire [15:0] _GEN_262;
  wire [15:0] _GEN_263;
  wire [15:0] _GEN_264;
  wire [15:0] _GEN_265;
  wire [15:0] _GEN_266;
  wire [15:0] _GEN_267;
  wire [15:0] _GEN_268;
  wire [15:0] _GEN_269;
  wire [15:0] _GEN_270;
  wire [15:0] _GEN_271;
  wire [15:0] _GEN_272;
  wire [15:0] _GEN_273;
  wire [15:0] _GEN_274;
  wire [15:0] _GEN_275;
  wire [15:0] _GEN_276;
  wire [15:0] _GEN_277;
  wire [15:0] _GEN_278;
  wire [15:0] _GEN_279;
  wire [15:0] _GEN_280;
  wire [15:0] _GEN_281;
  wire [15:0] _GEN_282;
  wire [15:0] _GEN_283;
  wire [15:0] _GEN_284;
  wire [15:0] _GEN_285;
  wire [15:0] _GEN_286;
  wire [15:0] _GEN_287;
  wire [15:0] _GEN_288;
  wire [15:0] _GEN_289;
  wire [15:0] _GEN_290;
  wire [15:0] _GEN_291;
  wire [15:0] _GEN_292;
  wire [15:0] _GEN_293;
  wire [15:0] _GEN_294;
  wire [15:0] _GEN_295;
  wire [15:0] _GEN_296;
  wire [15:0] _GEN_297;
  wire [15:0] _GEN_298;
  wire [15:0] _GEN_299;
  wire [15:0] _GEN_300;
  wire [15:0] _GEN_301;
  wire [15:0] _GEN_302;
  wire [15:0] _GEN_303;
  wire [15:0] _GEN_304;
  wire [15:0] _GEN_305;
  wire [15:0] _GEN_306;
  wire [15:0] _GEN_307;
  wire [15:0] _GEN_308;
  wire [15:0] _GEN_309;
  wire [15:0] _GEN_310;
  wire [15:0] _GEN_311;
  wire [15:0] _GEN_312;
  wire [15:0] _GEN_313;
  wire [15:0] _GEN_314;
  wire [15:0] _GEN_315;
  wire [15:0] _GEN_316;
  wire [15:0] _GEN_317;
  wire [15:0] _GEN_318;
  wire [15:0] _GEN_319;
  wire [15:0] _GEN_320;
  wire [15:0] _GEN_321;
  wire [15:0] _GEN_322;
  wire [15:0] _GEN_323;
  wire [15:0] _GEN_324;
  wire [15:0] _GEN_325;
  wire [15:0] _GEN_326;
  wire [15:0] _GEN_327;
  wire [15:0] _GEN_328;
  wire [15:0] _GEN_329;
  wire [15:0] _GEN_330;
  wire [15:0] _GEN_331;
  wire [15:0] _GEN_332;
  wire [15:0] _GEN_333;
  wire [15:0] _GEN_334;
  wire [15:0] _GEN_335;
  wire [15:0] _GEN_336;
  wire [15:0] _GEN_337;
  wire [15:0] _GEN_338;
  wire [15:0] _GEN_339;
  wire [15:0] _GEN_340;
  wire [15:0] _GEN_341;
  wire [15:0] _GEN_342;
  wire [15:0] _GEN_343;
  wire [15:0] _GEN_344;
  wire [15:0] _GEN_345;
  wire [15:0] _GEN_346;
  wire [15:0] _GEN_347;
  wire [15:0] _GEN_348;
  wire [15:0] _GEN_349;
  wire [15:0] _GEN_350;
  wire [15:0] _GEN_351;
  wire [15:0] _GEN_352;
  wire [15:0] _GEN_353;
  wire [15:0] _GEN_354;
  wire [15:0] _GEN_355;
  wire [15:0] _GEN_356;
  wire [15:0] _GEN_357;
  wire [15:0] _GEN_358;
  wire [15:0] _GEN_359;
  wire [15:0] _GEN_360;
  wire [15:0] _GEN_361;
  wire [15:0] _GEN_362;
  wire [15:0] _GEN_363;
  wire [15:0] _GEN_364;
  wire [15:0] _GEN_365;
  wire [15:0] _GEN_366;
  wire [15:0] _GEN_367;
  wire [15:0] _GEN_368;
  wire [15:0] _GEN_369;
  wire [15:0] _GEN_370;
  wire [15:0] _GEN_371;
  wire [15:0] _GEN_372;
  wire [15:0] _GEN_373;
  wire [15:0] _GEN_374;
  wire [15:0] _GEN_375;
  wire [15:0] _GEN_376;
  wire [15:0] _GEN_377;
  wire [15:0] _GEN_378;
  wire [15:0] _GEN_379;
  wire [15:0] _GEN_380;
  wire [15:0] _GEN_381;
  wire [15:0] _GEN_382;
  wire [15:0] _GEN_383;
  wire [15:0] _GEN_384;
  wire [15:0] _GEN_385;
  wire [15:0] _GEN_386;
  wire [15:0] _GEN_387;
  wire [15:0] _GEN_388;
  wire [15:0] _GEN_389;
  wire [15:0] _GEN_390;
  wire [15:0] _GEN_391;
  wire [15:0] _GEN_392;
  wire [15:0] _GEN_393;
  wire [15:0] _GEN_394;
  wire [15:0] _GEN_395;
  wire [15:0] _GEN_396;
  wire [15:0] _GEN_397;
  wire [15:0] _GEN_398;
  wire [15:0] _GEN_399;
  wire [15:0] _GEN_401;
  wire [15:0] _GEN_402;
  wire [15:0] _GEN_403;
  wire [15:0] _GEN_404;
  wire [15:0] _GEN_405;
  wire [15:0] _GEN_406;
  wire [15:0] _GEN_407;
  wire [15:0] _GEN_408;
  wire [15:0] _GEN_409;
  wire [15:0] _GEN_410;
  wire [15:0] _GEN_411;
  wire [15:0] _GEN_412;
  wire [15:0] _GEN_413;
  wire [15:0] _GEN_414;
  wire [15:0] _GEN_415;
  wire [15:0] _GEN_416;
  wire [15:0] _GEN_417;
  wire [15:0] _GEN_418;
  wire [15:0] _GEN_419;
  wire [15:0] _GEN_420;
  wire [15:0] _GEN_421;
  wire [15:0] _GEN_422;
  wire [15:0] _GEN_423;
  wire [15:0] _GEN_424;
  wire [15:0] _GEN_425;
  wire [15:0] _GEN_426;
  wire [15:0] _GEN_427;
  wire [15:0] _GEN_428;
  wire [15:0] _GEN_429;
  wire [15:0] _GEN_430;
  wire [15:0] _GEN_431;
  wire [15:0] _GEN_432;
  wire [15:0] _GEN_433;
  wire [15:0] _GEN_434;
  wire [15:0] _GEN_435;
  wire [15:0] _GEN_436;
  wire [15:0] _GEN_437;
  wire [15:0] _GEN_438;
  wire [15:0] _GEN_439;
  wire [15:0] _GEN_440;
  wire [15:0] _GEN_441;
  wire [15:0] _GEN_442;
  wire [15:0] _GEN_443;
  wire [15:0] _GEN_444;
  wire [15:0] _GEN_445;
  wire [15:0] _GEN_446;
  wire [15:0] _GEN_447;
  wire [15:0] _GEN_448;
  wire [15:0] _GEN_449;
  wire [15:0] _GEN_450;
  wire [15:0] _GEN_451;
  wire [15:0] _GEN_452;
  wire [15:0] _GEN_453;
  wire [15:0] _GEN_454;
  wire [15:0] _GEN_455;
  wire [15:0] _GEN_456;
  wire [15:0] _GEN_457;
  wire [15:0] _GEN_458;
  wire [15:0] _GEN_459;
  wire [15:0] _GEN_460;
  wire [15:0] _GEN_461;
  wire [15:0] _GEN_462;
  wire [15:0] _GEN_463;
  wire [15:0] _GEN_464;
  wire [15:0] _GEN_465;
  wire [15:0] _GEN_466;
  wire [15:0] _GEN_467;
  wire [15:0] _GEN_468;
  wire [15:0] _GEN_469;
  wire [15:0] _GEN_470;
  wire [15:0] _GEN_471;
  wire [15:0] _GEN_472;
  wire [15:0] _GEN_473;
  wire [15:0] _GEN_474;
  wire [15:0] _GEN_475;
  wire [15:0] _GEN_476;
  wire [15:0] _GEN_477;
  wire [15:0] _GEN_478;
  wire [15:0] _GEN_479;
  wire [15:0] _GEN_480;
  wire [15:0] _GEN_481;
  wire [15:0] _GEN_482;
  wire [15:0] _GEN_483;
  wire [15:0] _GEN_484;
  wire [15:0] _GEN_485;
  wire [15:0] _GEN_486;
  wire [15:0] _GEN_487;
  wire [15:0] _GEN_488;
  wire [15:0] _GEN_489;
  wire [15:0] _GEN_490;
  wire [15:0] _GEN_491;
  wire [15:0] _GEN_492;
  wire [15:0] _GEN_493;
  wire [15:0] _GEN_494;
  wire [15:0] _GEN_495;
  wire [15:0] _GEN_496;
  wire [15:0] _GEN_497;
  wire [15:0] _GEN_498;
  wire [15:0] _GEN_499;
  wire [15:0] _GEN_500;
  wire [15:0] _GEN_501;
  wire [15:0] _GEN_502;
  wire [15:0] _GEN_503;
  wire [15:0] _GEN_504;
  wire [15:0] _GEN_505;
  wire [15:0] _GEN_506;
  wire [15:0] _GEN_507;
  wire [15:0] _GEN_508;
  wire [15:0] _GEN_509;
  wire [15:0] _GEN_510;
  wire [15:0] _GEN_511;
  wire [15:0] _GEN_512;
  wire [15:0] _GEN_513;
  wire [15:0] _GEN_514;
  wire [15:0] _GEN_515;
  wire [15:0] _GEN_516;
  wire [15:0] _GEN_517;
  wire [15:0] _GEN_518;
  wire [15:0] _GEN_519;
  wire [15:0] _GEN_520;
  wire [15:0] _GEN_521;
  wire [15:0] _GEN_522;
  wire [15:0] _GEN_523;
  wire [15:0] _GEN_524;
  wire [15:0] _GEN_525;
  wire [15:0] _GEN_526;
  wire [15:0] _GEN_527;
  wire [15:0] _GEN_528;
  wire [15:0] _GEN_529;
  wire [15:0] _GEN_530;
  wire [15:0] _GEN_531;
  wire [15:0] _GEN_532;
  wire [15:0] _GEN_533;
  wire [15:0] _GEN_534;
  wire [15:0] _GEN_535;
  wire [15:0] _GEN_536;
  wire [15:0] _GEN_537;
  wire [15:0] _GEN_538;
  wire [15:0] _GEN_539;
  wire [15:0] _GEN_540;
  wire [15:0] _GEN_541;
  wire [15:0] _GEN_542;
  wire [15:0] _GEN_543;
  wire [15:0] _GEN_544;
  wire [15:0] _GEN_545;
  wire [15:0] _GEN_546;
  wire [15:0] _GEN_547;
  wire [15:0] _GEN_548;
  wire [15:0] _GEN_549;
  wire [15:0] _GEN_550;
  wire [15:0] _GEN_551;
  wire [15:0] _GEN_552;
  wire [15:0] _GEN_553;
  wire [15:0] _GEN_554;
  wire [15:0] _GEN_555;
  wire [15:0] _GEN_556;
  wire [15:0] _GEN_557;
  wire [15:0] _GEN_558;
  wire [15:0] _GEN_559;
  wire [15:0] _GEN_560;
  wire [15:0] _GEN_561;
  wire [15:0] _GEN_562;
  wire [15:0] _GEN_563;
  wire [15:0] _GEN_564;
  wire [15:0] _GEN_565;
  wire [15:0] _GEN_566;
  wire [15:0] _GEN_567;
  wire [15:0] _GEN_568;
  wire [15:0] _GEN_569;
  wire [15:0] _GEN_570;
  wire [15:0] _GEN_571;
  wire [15:0] _GEN_572;
  wire [15:0] _GEN_573;
  wire [15:0] _GEN_574;
  wire [15:0] _GEN_575;
  wire [15:0] _GEN_576;
  wire [15:0] _GEN_577;
  wire [15:0] _GEN_578;
  wire [15:0] _GEN_579;
  wire [15:0] _GEN_580;
  wire [15:0] _GEN_581;
  wire [15:0] _GEN_582;
  wire [15:0] _GEN_583;
  wire [15:0] _GEN_584;
  wire [15:0] _GEN_585;
  wire [15:0] _GEN_586;
  wire [15:0] _GEN_587;
  wire [15:0] _GEN_588;
  wire [15:0] _GEN_589;
  wire [15:0] _GEN_590;
  wire [15:0] _GEN_591;
  wire [15:0] _GEN_592;
  wire [15:0] _GEN_593;
  wire [15:0] _GEN_594;
  wire [15:0] _GEN_595;
  wire [15:0] _GEN_596;
  wire [15:0] _GEN_597;
  wire [15:0] _GEN_598;
  wire [15:0] _GEN_599;
  wire [15:0] _GEN_600;
  wire [15:0] _GEN_601;
  wire [15:0] _GEN_602;
  wire [15:0] _GEN_603;
  wire [15:0] _GEN_604;
  wire [15:0] _GEN_605;
  wire [15:0] _GEN_606;
  wire [15:0] _GEN_607;
  wire [15:0] _GEN_608;
  wire [15:0] _GEN_609;
  wire [15:0] _GEN_610;
  wire [15:0] _GEN_611;
  wire [15:0] _GEN_612;
  wire [15:0] _GEN_613;
  wire [15:0] _GEN_614;
  wire [15:0] _GEN_615;
  wire [15:0] _GEN_616;
  wire [15:0] _GEN_617;
  wire [15:0] _GEN_618;
  wire [15:0] _GEN_619;
  wire [15:0] _GEN_620;
  wire [15:0] _GEN_621;
  wire [15:0] _GEN_622;
  wire [15:0] _GEN_623;
  wire [15:0] _GEN_624;
  wire [15:0] _GEN_625;
  wire [15:0] _GEN_626;
  wire [15:0] _GEN_627;
  wire [15:0] _GEN_628;
  wire [15:0] _GEN_629;
  wire [15:0] _GEN_630;
  wire [15:0] _GEN_631;
  wire [15:0] _GEN_632;
  wire [15:0] _GEN_633;
  wire [15:0] _GEN_634;
  wire [15:0] _GEN_635;
  wire [15:0] _GEN_636;
  wire [15:0] _GEN_637;
  wire [15:0] _GEN_638;
  wire [15:0] _GEN_639;
  wire [15:0] _GEN_640;
  wire [15:0] _GEN_641;
  wire [15:0] _GEN_642;
  wire [15:0] _GEN_643;
  wire [15:0] _GEN_644;
  wire [15:0] _GEN_645;
  wire [15:0] _GEN_646;
  wire [15:0] _GEN_647;
  wire [15:0] _GEN_648;
  wire [15:0] _GEN_649;
  wire [15:0] _GEN_650;
  wire [15:0] _GEN_651;
  wire [15:0] _GEN_652;
  wire [15:0] _GEN_653;
  wire [15:0] _GEN_654;
  wire [15:0] _GEN_655;
  wire [15:0] _GEN_656;
  wire [15:0] _GEN_657;
  wire [15:0] _GEN_658;
  wire [15:0] _GEN_659;
  wire [15:0] _GEN_660;
  wire [15:0] _GEN_661;
  wire [15:0] _GEN_662;
  wire [15:0] _GEN_663;
  wire [15:0] _GEN_664;
  wire [15:0] _GEN_665;
  wire [15:0] _GEN_666;
  wire [15:0] _GEN_667;
  wire [15:0] _GEN_668;
  wire [15:0] _GEN_669;
  wire [15:0] _GEN_670;
  wire [15:0] _GEN_671;
  wire [15:0] _GEN_672;
  wire [15:0] _GEN_673;
  wire [15:0] _GEN_674;
  wire [15:0] _GEN_675;
  wire [15:0] _GEN_676;
  wire [15:0] _GEN_677;
  wire [15:0] _GEN_678;
  wire [15:0] _GEN_679;
  wire [15:0] _GEN_680;
  wire [15:0] _GEN_681;
  wire [15:0] _GEN_682;
  wire [15:0] _GEN_683;
  wire [15:0] _GEN_684;
  wire [15:0] _GEN_685;
  wire [15:0] _GEN_686;
  wire [15:0] _GEN_687;
  wire [15:0] _GEN_688;
  wire [15:0] _GEN_689;
  wire [15:0] _GEN_690;
  wire [15:0] _GEN_691;
  wire [15:0] _GEN_692;
  wire [15:0] _GEN_693;
  wire [15:0] _GEN_694;
  wire [15:0] _GEN_695;
  wire [15:0] _GEN_696;
  wire [15:0] _GEN_697;
  wire [15:0] _GEN_698;
  wire [15:0] _GEN_699;
  wire [15:0] _GEN_700;
  wire [15:0] _GEN_701;
  wire [15:0] _GEN_702;
  wire [15:0] _GEN_703;
  wire [15:0] _GEN_704;
  wire [15:0] _GEN_705;
  wire [15:0] _GEN_706;
  wire [15:0] _GEN_707;
  wire [15:0] _GEN_708;
  wire [15:0] _GEN_709;
  wire [15:0] _GEN_710;
  wire [15:0] _GEN_711;
  wire [15:0] _GEN_712;
  wire [15:0] _GEN_713;
  wire [15:0] _GEN_714;
  wire [15:0] _GEN_715;
  wire [15:0] _GEN_716;
  wire [15:0] _GEN_717;
  wire [15:0] _GEN_718;
  wire [15:0] _GEN_719;
  wire [15:0] _GEN_720;
  wire [15:0] _GEN_721;
  wire [15:0] _GEN_722;
  wire [15:0] _GEN_723;
  wire [15:0] _GEN_724;
  wire [15:0] _GEN_725;
  wire [15:0] _GEN_726;
  wire [15:0] _GEN_727;
  wire [15:0] _GEN_728;
  wire [15:0] _GEN_729;
  wire [15:0] _GEN_730;
  wire [15:0] _GEN_731;
  wire [15:0] _GEN_732;
  wire [15:0] _GEN_733;
  wire [15:0] _GEN_734;
  wire [15:0] _GEN_735;
  wire [15:0] _GEN_736;
  wire [15:0] _GEN_737;
  wire [15:0] _GEN_738;
  wire [15:0] _GEN_739;
  wire [15:0] _GEN_740;
  wire [15:0] _GEN_741;
  wire [15:0] _GEN_742;
  wire [15:0] _GEN_743;
  wire [15:0] _GEN_744;
  wire [15:0] _GEN_745;
  wire [15:0] _GEN_746;
  wire [15:0] _GEN_747;
  wire [15:0] _GEN_748;
  wire [15:0] _GEN_749;
  wire [15:0] _GEN_750;
  wire [15:0] _GEN_751;
  wire [15:0] _GEN_752;
  wire [15:0] _GEN_753;
  wire [15:0] _GEN_754;
  wire [15:0] _GEN_755;
  wire [15:0] _GEN_756;
  wire [15:0] _GEN_757;
  wire [15:0] _GEN_758;
  wire [15:0] _GEN_759;
  wire [15:0] _GEN_760;
  wire [15:0] _GEN_761;
  wire [15:0] _GEN_762;
  wire [15:0] _GEN_763;
  wire [15:0] _GEN_764;
  wire [15:0] _GEN_765;
  wire [15:0] _GEN_766;
  wire [15:0] _GEN_767;
  wire [15:0] _GEN_768;
  wire [15:0] _GEN_769;
  wire [15:0] _GEN_770;
  wire [15:0] _GEN_771;
  wire [15:0] _GEN_772;
  wire [15:0] _GEN_773;
  wire [15:0] _GEN_774;
  wire [15:0] _GEN_775;
  wire [15:0] _GEN_776;
  wire [15:0] _GEN_777;
  wire [15:0] _GEN_778;
  wire [15:0] _GEN_779;
  wire [15:0] _GEN_780;
  wire [15:0] _GEN_781;
  wire [15:0] _GEN_782;
  wire [15:0] _GEN_783;
  wire [15:0] _GEN_784;
  wire [15:0] _GEN_785;
  wire [15:0] _GEN_786;
  wire [15:0] _GEN_787;
  wire [15:0] _GEN_788;
  wire [15:0] _GEN_789;
  wire [15:0] _GEN_790;
  wire [15:0] _GEN_791;
  wire [15:0] _GEN_792;
  wire [15:0] _GEN_793;
  wire [15:0] _GEN_794;
  wire [15:0] _GEN_795;
  wire [15:0] _GEN_796;
  wire [15:0] _GEN_797;
  wire [15:0] _GEN_798;
  wire [15:0] _GEN_799;
  wire [31:0] _T_800;
  wire [32:0] _T_801;
  wire [9:0] _T_802;
  wire [9:0] _GEN_800;
  wire [32:0] _GEN_801;
  wire [9:0] _GEN_802;
  wire [31:0] _GEN_804;
  wire [32:0] _GEN_805;
  wire [32:0] _GEN_806;
  wire [9:0] _GEN_807;
  assign a_0 = io_a[15:0];
  assign b_0 = io_b[15:0];
  assign a_1 = io_a[31:16];
  assign b_1 = io_b[31:16];
  assign a_2 = io_a[47:32];
  assign b_2 = io_b[47:32];
  assign a_3 = io_a[63:48];
  assign b_3 = io_b[63:48];
  assign a_4 = io_a[79:64];
  assign b_4 = io_b[79:64];
  assign a_5 = io_a[95:80];
  assign b_5 = io_b[95:80];
  assign a_6 = io_a[111:96];
  assign b_6 = io_b[111:96];
  assign a_7 = io_a[127:112];
  assign b_7 = io_b[127:112];
  assign a_8 = io_a[143:128];
  assign b_8 = io_b[143:128];
  assign a_9 = io_a[159:144];
  assign b_9 = io_b[159:144];
  assign a_10 = io_a[175:160];
  assign b_10 = io_b[175:160];
  assign a_11 = io_a[191:176];
  assign b_11 = io_b[191:176];
  assign a_12 = io_a[207:192];
  assign b_12 = io_b[207:192];
  assign a_13 = io_a[223:208];
  assign b_13 = io_b[223:208];
  assign a_14 = io_a[239:224];
  assign b_14 = io_b[239:224];
  assign a_15 = io_a[255:240];
  assign b_15 = io_b[255:240];
  assign a_16 = io_a[271:256];
  assign b_16 = io_b[271:256];
  assign a_17 = io_a[287:272];
  assign b_17 = io_b[287:272];
  assign a_18 = io_a[303:288];
  assign b_18 = io_b[303:288];
  assign a_19 = io_a[319:304];
  assign b_19 = io_b[319:304];
  assign a_20 = io_a[335:320];
  assign b_20 = io_b[335:320];
  assign a_21 = io_a[351:336];
  assign b_21 = io_b[351:336];
  assign a_22 = io_a[367:352];
  assign b_22 = io_b[367:352];
  assign a_23 = io_a[383:368];
  assign b_23 = io_b[383:368];
  assign a_24 = io_a[399:384];
  assign b_24 = io_b[399:384];
  assign a_25 = io_a[415:400];
  assign b_25 = io_b[415:400];
  assign a_26 = io_a[431:416];
  assign b_26 = io_b[431:416];
  assign a_27 = io_a[447:432];
  assign b_27 = io_b[447:432];
  assign a_28 = io_a[463:448];
  assign b_28 = io_b[463:448];
  assign a_29 = io_a[479:464];
  assign b_29 = io_b[479:464];
  assign a_30 = io_a[495:480];
  assign b_30 = io_b[495:480];
  assign a_31 = io_a[511:496];
  assign b_31 = io_b[511:496];
  assign a_32 = io_a[527:512];
  assign b_32 = io_b[527:512];
  assign a_33 = io_a[543:528];
  assign b_33 = io_b[543:528];
  assign a_34 = io_a[559:544];
  assign b_34 = io_b[559:544];
  assign a_35 = io_a[575:560];
  assign b_35 = io_b[575:560];
  assign a_36 = io_a[591:576];
  assign b_36 = io_b[591:576];
  assign a_37 = io_a[607:592];
  assign b_37 = io_b[607:592];
  assign a_38 = io_a[623:608];
  assign b_38 = io_b[623:608];
  assign a_39 = io_a[639:624];
  assign b_39 = io_b[639:624];
  assign a_40 = io_a[655:640];
  assign b_40 = io_b[655:640];
  assign a_41 = io_a[671:656];
  assign b_41 = io_b[671:656];
  assign a_42 = io_a[687:672];
  assign b_42 = io_b[687:672];
  assign a_43 = io_a[703:688];
  assign b_43 = io_b[703:688];
  assign a_44 = io_a[719:704];
  assign b_44 = io_b[719:704];
  assign a_45 = io_a[735:720];
  assign b_45 = io_b[735:720];
  assign a_46 = io_a[751:736];
  assign b_46 = io_b[751:736];
  assign a_47 = io_a[767:752];
  assign b_47 = io_b[767:752];
  assign a_48 = io_a[783:768];
  assign b_48 = io_b[783:768];
  assign a_49 = io_a[799:784];
  assign b_49 = io_b[799:784];
  assign a_50 = io_a[815:800];
  assign b_50 = io_b[815:800];
  assign a_51 = io_a[831:816];
  assign b_51 = io_b[831:816];
  assign a_52 = io_a[847:832];
  assign b_52 = io_b[847:832];
  assign a_53 = io_a[863:848];
  assign b_53 = io_b[863:848];
  assign a_54 = io_a[879:864];
  assign b_54 = io_b[879:864];
  assign a_55 = io_a[895:880];
  assign b_55 = io_b[895:880];
  assign a_56 = io_a[911:896];
  assign b_56 = io_b[911:896];
  assign a_57 = io_a[927:912];
  assign b_57 = io_b[927:912];
  assign a_58 = io_a[943:928];
  assign b_58 = io_b[943:928];
  assign a_59 = io_a[959:944];
  assign b_59 = io_b[959:944];
  assign a_60 = io_a[975:960];
  assign b_60 = io_b[975:960];
  assign a_61 = io_a[991:976];
  assign b_61 = io_b[991:976];
  assign a_62 = io_a[1007:992];
  assign b_62 = io_b[1007:992];
  assign a_63 = io_a[1023:1008];
  assign b_63 = io_b[1023:1008];
  assign a_64 = io_a[1039:1024];
  assign b_64 = io_b[1039:1024];
  assign a_65 = io_a[1055:1040];
  assign b_65 = io_b[1055:1040];
  assign a_66 = io_a[1071:1056];
  assign b_66 = io_b[1071:1056];
  assign a_67 = io_a[1087:1072];
  assign b_67 = io_b[1087:1072];
  assign a_68 = io_a[1103:1088];
  assign b_68 = io_b[1103:1088];
  assign a_69 = io_a[1119:1104];
  assign b_69 = io_b[1119:1104];
  assign a_70 = io_a[1135:1120];
  assign b_70 = io_b[1135:1120];
  assign a_71 = io_a[1151:1136];
  assign b_71 = io_b[1151:1136];
  assign a_72 = io_a[1167:1152];
  assign b_72 = io_b[1167:1152];
  assign a_73 = io_a[1183:1168];
  assign b_73 = io_b[1183:1168];
  assign a_74 = io_a[1199:1184];
  assign b_74 = io_b[1199:1184];
  assign a_75 = io_a[1215:1200];
  assign b_75 = io_b[1215:1200];
  assign a_76 = io_a[1231:1216];
  assign b_76 = io_b[1231:1216];
  assign a_77 = io_a[1247:1232];
  assign b_77 = io_b[1247:1232];
  assign a_78 = io_a[1263:1248];
  assign b_78 = io_b[1263:1248];
  assign a_79 = io_a[1279:1264];
  assign b_79 = io_b[1279:1264];
  assign a_80 = io_a[1295:1280];
  assign b_80 = io_b[1295:1280];
  assign a_81 = io_a[1311:1296];
  assign b_81 = io_b[1311:1296];
  assign a_82 = io_a[1327:1312];
  assign b_82 = io_b[1327:1312];
  assign a_83 = io_a[1343:1328];
  assign b_83 = io_b[1343:1328];
  assign a_84 = io_a[1359:1344];
  assign b_84 = io_b[1359:1344];
  assign a_85 = io_a[1375:1360];
  assign b_85 = io_b[1375:1360];
  assign a_86 = io_a[1391:1376];
  assign b_86 = io_b[1391:1376];
  assign a_87 = io_a[1407:1392];
  assign b_87 = io_b[1407:1392];
  assign a_88 = io_a[1423:1408];
  assign b_88 = io_b[1423:1408];
  assign a_89 = io_a[1439:1424];
  assign b_89 = io_b[1439:1424];
  assign a_90 = io_a[1455:1440];
  assign b_90 = io_b[1455:1440];
  assign a_91 = io_a[1471:1456];
  assign b_91 = io_b[1471:1456];
  assign a_92 = io_a[1487:1472];
  assign b_92 = io_b[1487:1472];
  assign a_93 = io_a[1503:1488];
  assign b_93 = io_b[1503:1488];
  assign a_94 = io_a[1519:1504];
  assign b_94 = io_b[1519:1504];
  assign a_95 = io_a[1535:1520];
  assign b_95 = io_b[1535:1520];
  assign a_96 = io_a[1551:1536];
  assign b_96 = io_b[1551:1536];
  assign a_97 = io_a[1567:1552];
  assign b_97 = io_b[1567:1552];
  assign a_98 = io_a[1583:1568];
  assign b_98 = io_b[1583:1568];
  assign a_99 = io_a[1599:1584];
  assign b_99 = io_b[1599:1584];
  assign a_100 = io_a[1615:1600];
  assign b_100 = io_b[1615:1600];
  assign a_101 = io_a[1631:1616];
  assign b_101 = io_b[1631:1616];
  assign a_102 = io_a[1647:1632];
  assign b_102 = io_b[1647:1632];
  assign a_103 = io_a[1663:1648];
  assign b_103 = io_b[1663:1648];
  assign a_104 = io_a[1679:1664];
  assign b_104 = io_b[1679:1664];
  assign a_105 = io_a[1695:1680];
  assign b_105 = io_b[1695:1680];
  assign a_106 = io_a[1711:1696];
  assign b_106 = io_b[1711:1696];
  assign a_107 = io_a[1727:1712];
  assign b_107 = io_b[1727:1712];
  assign a_108 = io_a[1743:1728];
  assign b_108 = io_b[1743:1728];
  assign a_109 = io_a[1759:1744];
  assign b_109 = io_b[1759:1744];
  assign a_110 = io_a[1775:1760];
  assign b_110 = io_b[1775:1760];
  assign a_111 = io_a[1791:1776];
  assign b_111 = io_b[1791:1776];
  assign a_112 = io_a[1807:1792];
  assign b_112 = io_b[1807:1792];
  assign a_113 = io_a[1823:1808];
  assign b_113 = io_b[1823:1808];
  assign a_114 = io_a[1839:1824];
  assign b_114 = io_b[1839:1824];
  assign a_115 = io_a[1855:1840];
  assign b_115 = io_b[1855:1840];
  assign a_116 = io_a[1871:1856];
  assign b_116 = io_b[1871:1856];
  assign a_117 = io_a[1887:1872];
  assign b_117 = io_b[1887:1872];
  assign a_118 = io_a[1903:1888];
  assign b_118 = io_b[1903:1888];
  assign a_119 = io_a[1919:1904];
  assign b_119 = io_b[1919:1904];
  assign a_120 = io_a[1935:1920];
  assign b_120 = io_b[1935:1920];
  assign a_121 = io_a[1951:1936];
  assign b_121 = io_b[1951:1936];
  assign a_122 = io_a[1967:1952];
  assign b_122 = io_b[1967:1952];
  assign a_123 = io_a[1983:1968];
  assign b_123 = io_b[1983:1968];
  assign a_124 = io_a[1999:1984];
  assign b_124 = io_b[1999:1984];
  assign a_125 = io_a[2015:2000];
  assign b_125 = io_b[2015:2000];
  assign a_126 = io_a[2031:2016];
  assign b_126 = io_b[2031:2016];
  assign a_127 = io_a[2047:2032];
  assign b_127 = io_b[2047:2032];
  assign a_128 = io_a[2063:2048];
  assign b_128 = io_b[2063:2048];
  assign a_129 = io_a[2079:2064];
  assign b_129 = io_b[2079:2064];
  assign a_130 = io_a[2095:2080];
  assign b_130 = io_b[2095:2080];
  assign a_131 = io_a[2111:2096];
  assign b_131 = io_b[2111:2096];
  assign a_132 = io_a[2127:2112];
  assign b_132 = io_b[2127:2112];
  assign a_133 = io_a[2143:2128];
  assign b_133 = io_b[2143:2128];
  assign a_134 = io_a[2159:2144];
  assign b_134 = io_b[2159:2144];
  assign a_135 = io_a[2175:2160];
  assign b_135 = io_b[2175:2160];
  assign a_136 = io_a[2191:2176];
  assign b_136 = io_b[2191:2176];
  assign a_137 = io_a[2207:2192];
  assign b_137 = io_b[2207:2192];
  assign a_138 = io_a[2223:2208];
  assign b_138 = io_b[2223:2208];
  assign a_139 = io_a[2239:2224];
  assign b_139 = io_b[2239:2224];
  assign a_140 = io_a[2255:2240];
  assign b_140 = io_b[2255:2240];
  assign a_141 = io_a[2271:2256];
  assign b_141 = io_b[2271:2256];
  assign a_142 = io_a[2287:2272];
  assign b_142 = io_b[2287:2272];
  assign a_143 = io_a[2303:2288];
  assign b_143 = io_b[2303:2288];
  assign a_144 = io_a[2319:2304];
  assign b_144 = io_b[2319:2304];
  assign a_145 = io_a[2335:2320];
  assign b_145 = io_b[2335:2320];
  assign a_146 = io_a[2351:2336];
  assign b_146 = io_b[2351:2336];
  assign a_147 = io_a[2367:2352];
  assign b_147 = io_b[2367:2352];
  assign a_148 = io_a[2383:2368];
  assign b_148 = io_b[2383:2368];
  assign a_149 = io_a[2399:2384];
  assign b_149 = io_b[2399:2384];
  assign a_150 = io_a[2415:2400];
  assign b_150 = io_b[2415:2400];
  assign a_151 = io_a[2431:2416];
  assign b_151 = io_b[2431:2416];
  assign a_152 = io_a[2447:2432];
  assign b_152 = io_b[2447:2432];
  assign a_153 = io_a[2463:2448];
  assign b_153 = io_b[2463:2448];
  assign a_154 = io_a[2479:2464];
  assign b_154 = io_b[2479:2464];
  assign a_155 = io_a[2495:2480];
  assign b_155 = io_b[2495:2480];
  assign a_156 = io_a[2511:2496];
  assign b_156 = io_b[2511:2496];
  assign a_157 = io_a[2527:2512];
  assign b_157 = io_b[2527:2512];
  assign a_158 = io_a[2543:2528];
  assign b_158 = io_b[2543:2528];
  assign a_159 = io_a[2559:2544];
  assign b_159 = io_b[2559:2544];
  assign a_160 = io_a[2575:2560];
  assign b_160 = io_b[2575:2560];
  assign a_161 = io_a[2591:2576];
  assign b_161 = io_b[2591:2576];
  assign a_162 = io_a[2607:2592];
  assign b_162 = io_b[2607:2592];
  assign a_163 = io_a[2623:2608];
  assign b_163 = io_b[2623:2608];
  assign a_164 = io_a[2639:2624];
  assign b_164 = io_b[2639:2624];
  assign a_165 = io_a[2655:2640];
  assign b_165 = io_b[2655:2640];
  assign a_166 = io_a[2671:2656];
  assign b_166 = io_b[2671:2656];
  assign a_167 = io_a[2687:2672];
  assign b_167 = io_b[2687:2672];
  assign a_168 = io_a[2703:2688];
  assign b_168 = io_b[2703:2688];
  assign a_169 = io_a[2719:2704];
  assign b_169 = io_b[2719:2704];
  assign a_170 = io_a[2735:2720];
  assign b_170 = io_b[2735:2720];
  assign a_171 = io_a[2751:2736];
  assign b_171 = io_b[2751:2736];
  assign a_172 = io_a[2767:2752];
  assign b_172 = io_b[2767:2752];
  assign a_173 = io_a[2783:2768];
  assign b_173 = io_b[2783:2768];
  assign a_174 = io_a[2799:2784];
  assign b_174 = io_b[2799:2784];
  assign a_175 = io_a[2815:2800];
  assign b_175 = io_b[2815:2800];
  assign a_176 = io_a[2831:2816];
  assign b_176 = io_b[2831:2816];
  assign a_177 = io_a[2847:2832];
  assign b_177 = io_b[2847:2832];
  assign a_178 = io_a[2863:2848];
  assign b_178 = io_b[2863:2848];
  assign a_179 = io_a[2879:2864];
  assign b_179 = io_b[2879:2864];
  assign a_180 = io_a[2895:2880];
  assign b_180 = io_b[2895:2880];
  assign a_181 = io_a[2911:2896];
  assign b_181 = io_b[2911:2896];
  assign a_182 = io_a[2927:2912];
  assign b_182 = io_b[2927:2912];
  assign a_183 = io_a[2943:2928];
  assign b_183 = io_b[2943:2928];
  assign a_184 = io_a[2959:2944];
  assign b_184 = io_b[2959:2944];
  assign a_185 = io_a[2975:2960];
  assign b_185 = io_b[2975:2960];
  assign a_186 = io_a[2991:2976];
  assign b_186 = io_b[2991:2976];
  assign a_187 = io_a[3007:2992];
  assign b_187 = io_b[3007:2992];
  assign a_188 = io_a[3023:3008];
  assign b_188 = io_b[3023:3008];
  assign a_189 = io_a[3039:3024];
  assign b_189 = io_b[3039:3024];
  assign a_190 = io_a[3055:3040];
  assign b_190 = io_b[3055:3040];
  assign a_191 = io_a[3071:3056];
  assign b_191 = io_b[3071:3056];
  assign a_192 = io_a[3087:3072];
  assign b_192 = io_b[3087:3072];
  assign a_193 = io_a[3103:3088];
  assign b_193 = io_b[3103:3088];
  assign a_194 = io_a[3119:3104];
  assign b_194 = io_b[3119:3104];
  assign a_195 = io_a[3135:3120];
  assign b_195 = io_b[3135:3120];
  assign a_196 = io_a[3151:3136];
  assign b_196 = io_b[3151:3136];
  assign a_197 = io_a[3167:3152];
  assign b_197 = io_b[3167:3152];
  assign a_198 = io_a[3183:3168];
  assign b_198 = io_b[3183:3168];
  assign a_199 = io_a[3199:3184];
  assign b_199 = io_b[3199:3184];
  assign a_200 = io_a[3215:3200];
  assign b_200 = io_b[3215:3200];
  assign a_201 = io_a[3231:3216];
  assign b_201 = io_b[3231:3216];
  assign a_202 = io_a[3247:3232];
  assign b_202 = io_b[3247:3232];
  assign a_203 = io_a[3263:3248];
  assign b_203 = io_b[3263:3248];
  assign a_204 = io_a[3279:3264];
  assign b_204 = io_b[3279:3264];
  assign a_205 = io_a[3295:3280];
  assign b_205 = io_b[3295:3280];
  assign a_206 = io_a[3311:3296];
  assign b_206 = io_b[3311:3296];
  assign a_207 = io_a[3327:3312];
  assign b_207 = io_b[3327:3312];
  assign a_208 = io_a[3343:3328];
  assign b_208 = io_b[3343:3328];
  assign a_209 = io_a[3359:3344];
  assign b_209 = io_b[3359:3344];
  assign a_210 = io_a[3375:3360];
  assign b_210 = io_b[3375:3360];
  assign a_211 = io_a[3391:3376];
  assign b_211 = io_b[3391:3376];
  assign a_212 = io_a[3407:3392];
  assign b_212 = io_b[3407:3392];
  assign a_213 = io_a[3423:3408];
  assign b_213 = io_b[3423:3408];
  assign a_214 = io_a[3439:3424];
  assign b_214 = io_b[3439:3424];
  assign a_215 = io_a[3455:3440];
  assign b_215 = io_b[3455:3440];
  assign a_216 = io_a[3471:3456];
  assign b_216 = io_b[3471:3456];
  assign a_217 = io_a[3487:3472];
  assign b_217 = io_b[3487:3472];
  assign a_218 = io_a[3503:3488];
  assign b_218 = io_b[3503:3488];
  assign a_219 = io_a[3519:3504];
  assign b_219 = io_b[3519:3504];
  assign a_220 = io_a[3535:3520];
  assign b_220 = io_b[3535:3520];
  assign a_221 = io_a[3551:3536];
  assign b_221 = io_b[3551:3536];
  assign a_222 = io_a[3567:3552];
  assign b_222 = io_b[3567:3552];
  assign a_223 = io_a[3583:3568];
  assign b_223 = io_b[3583:3568];
  assign a_224 = io_a[3599:3584];
  assign b_224 = io_b[3599:3584];
  assign a_225 = io_a[3615:3600];
  assign b_225 = io_b[3615:3600];
  assign a_226 = io_a[3631:3616];
  assign b_226 = io_b[3631:3616];
  assign a_227 = io_a[3647:3632];
  assign b_227 = io_b[3647:3632];
  assign a_228 = io_a[3663:3648];
  assign b_228 = io_b[3663:3648];
  assign a_229 = io_a[3679:3664];
  assign b_229 = io_b[3679:3664];
  assign a_230 = io_a[3695:3680];
  assign b_230 = io_b[3695:3680];
  assign a_231 = io_a[3711:3696];
  assign b_231 = io_b[3711:3696];
  assign a_232 = io_a[3727:3712];
  assign b_232 = io_b[3727:3712];
  assign a_233 = io_a[3743:3728];
  assign b_233 = io_b[3743:3728];
  assign a_234 = io_a[3759:3744];
  assign b_234 = io_b[3759:3744];
  assign a_235 = io_a[3775:3760];
  assign b_235 = io_b[3775:3760];
  assign a_236 = io_a[3791:3776];
  assign b_236 = io_b[3791:3776];
  assign a_237 = io_a[3807:3792];
  assign b_237 = io_b[3807:3792];
  assign a_238 = io_a[3823:3808];
  assign b_238 = io_b[3823:3808];
  assign a_239 = io_a[3839:3824];
  assign b_239 = io_b[3839:3824];
  assign a_240 = io_a[3855:3840];
  assign b_240 = io_b[3855:3840];
  assign a_241 = io_a[3871:3856];
  assign b_241 = io_b[3871:3856];
  assign a_242 = io_a[3887:3872];
  assign b_242 = io_b[3887:3872];
  assign a_243 = io_a[3903:3888];
  assign b_243 = io_b[3903:3888];
  assign a_244 = io_a[3919:3904];
  assign b_244 = io_b[3919:3904];
  assign a_245 = io_a[3935:3920];
  assign b_245 = io_b[3935:3920];
  assign a_246 = io_a[3951:3936];
  assign b_246 = io_b[3951:3936];
  assign a_247 = io_a[3967:3952];
  assign b_247 = io_b[3967:3952];
  assign a_248 = io_a[3983:3968];
  assign b_248 = io_b[3983:3968];
  assign a_249 = io_a[3999:3984];
  assign b_249 = io_b[3999:3984];
  assign a_250 = io_a[4015:4000];
  assign b_250 = io_b[4015:4000];
  assign a_251 = io_a[4031:4016];
  assign b_251 = io_b[4031:4016];
  assign a_252 = io_a[4047:4032];
  assign b_252 = io_b[4047:4032];
  assign a_253 = io_a[4063:4048];
  assign b_253 = io_b[4063:4048];
  assign a_254 = io_a[4079:4064];
  assign b_254 = io_b[4079:4064];
  assign a_255 = io_a[4095:4080];
  assign b_255 = io_b[4095:4080];
  assign a_256 = io_a[4111:4096];
  assign b_256 = io_b[4111:4096];
  assign a_257 = io_a[4127:4112];
  assign b_257 = io_b[4127:4112];
  assign a_258 = io_a[4143:4128];
  assign b_258 = io_b[4143:4128];
  assign a_259 = io_a[4159:4144];
  assign b_259 = io_b[4159:4144];
  assign a_260 = io_a[4175:4160];
  assign b_260 = io_b[4175:4160];
  assign a_261 = io_a[4191:4176];
  assign b_261 = io_b[4191:4176];
  assign a_262 = io_a[4207:4192];
  assign b_262 = io_b[4207:4192];
  assign a_263 = io_a[4223:4208];
  assign b_263 = io_b[4223:4208];
  assign a_264 = io_a[4239:4224];
  assign b_264 = io_b[4239:4224];
  assign a_265 = io_a[4255:4240];
  assign b_265 = io_b[4255:4240];
  assign a_266 = io_a[4271:4256];
  assign b_266 = io_b[4271:4256];
  assign a_267 = io_a[4287:4272];
  assign b_267 = io_b[4287:4272];
  assign a_268 = io_a[4303:4288];
  assign b_268 = io_b[4303:4288];
  assign a_269 = io_a[4319:4304];
  assign b_269 = io_b[4319:4304];
  assign a_270 = io_a[4335:4320];
  assign b_270 = io_b[4335:4320];
  assign a_271 = io_a[4351:4336];
  assign b_271 = io_b[4351:4336];
  assign a_272 = io_a[4367:4352];
  assign b_272 = io_b[4367:4352];
  assign a_273 = io_a[4383:4368];
  assign b_273 = io_b[4383:4368];
  assign a_274 = io_a[4399:4384];
  assign b_274 = io_b[4399:4384];
  assign a_275 = io_a[4415:4400];
  assign b_275 = io_b[4415:4400];
  assign a_276 = io_a[4431:4416];
  assign b_276 = io_b[4431:4416];
  assign a_277 = io_a[4447:4432];
  assign b_277 = io_b[4447:4432];
  assign a_278 = io_a[4463:4448];
  assign b_278 = io_b[4463:4448];
  assign a_279 = io_a[4479:4464];
  assign b_279 = io_b[4479:4464];
  assign a_280 = io_a[4495:4480];
  assign b_280 = io_b[4495:4480];
  assign a_281 = io_a[4511:4496];
  assign b_281 = io_b[4511:4496];
  assign a_282 = io_a[4527:4512];
  assign b_282 = io_b[4527:4512];
  assign a_283 = io_a[4543:4528];
  assign b_283 = io_b[4543:4528];
  assign a_284 = io_a[4559:4544];
  assign b_284 = io_b[4559:4544];
  assign a_285 = io_a[4575:4560];
  assign b_285 = io_b[4575:4560];
  assign a_286 = io_a[4591:4576];
  assign b_286 = io_b[4591:4576];
  assign a_287 = io_a[4607:4592];
  assign b_287 = io_b[4607:4592];
  assign a_288 = io_a[4623:4608];
  assign b_288 = io_b[4623:4608];
  assign a_289 = io_a[4639:4624];
  assign b_289 = io_b[4639:4624];
  assign a_290 = io_a[4655:4640];
  assign b_290 = io_b[4655:4640];
  assign a_291 = io_a[4671:4656];
  assign b_291 = io_b[4671:4656];
  assign a_292 = io_a[4687:4672];
  assign b_292 = io_b[4687:4672];
  assign a_293 = io_a[4703:4688];
  assign b_293 = io_b[4703:4688];
  assign a_294 = io_a[4719:4704];
  assign b_294 = io_b[4719:4704];
  assign a_295 = io_a[4735:4720];
  assign b_295 = io_b[4735:4720];
  assign a_296 = io_a[4751:4736];
  assign b_296 = io_b[4751:4736];
  assign a_297 = io_a[4767:4752];
  assign b_297 = io_b[4767:4752];
  assign a_298 = io_a[4783:4768];
  assign b_298 = io_b[4783:4768];
  assign a_299 = io_a[4799:4784];
  assign b_299 = io_b[4799:4784];
  assign a_300 = io_a[4815:4800];
  assign b_300 = io_b[4815:4800];
  assign a_301 = io_a[4831:4816];
  assign b_301 = io_b[4831:4816];
  assign a_302 = io_a[4847:4832];
  assign b_302 = io_b[4847:4832];
  assign a_303 = io_a[4863:4848];
  assign b_303 = io_b[4863:4848];
  assign a_304 = io_a[4879:4864];
  assign b_304 = io_b[4879:4864];
  assign a_305 = io_a[4895:4880];
  assign b_305 = io_b[4895:4880];
  assign a_306 = io_a[4911:4896];
  assign b_306 = io_b[4911:4896];
  assign a_307 = io_a[4927:4912];
  assign b_307 = io_b[4927:4912];
  assign a_308 = io_a[4943:4928];
  assign b_308 = io_b[4943:4928];
  assign a_309 = io_a[4959:4944];
  assign b_309 = io_b[4959:4944];
  assign a_310 = io_a[4975:4960];
  assign b_310 = io_b[4975:4960];
  assign a_311 = io_a[4991:4976];
  assign b_311 = io_b[4991:4976];
  assign a_312 = io_a[5007:4992];
  assign b_312 = io_b[5007:4992];
  assign a_313 = io_a[5023:5008];
  assign b_313 = io_b[5023:5008];
  assign a_314 = io_a[5039:5024];
  assign b_314 = io_b[5039:5024];
  assign a_315 = io_a[5055:5040];
  assign b_315 = io_b[5055:5040];
  assign a_316 = io_a[5071:5056];
  assign b_316 = io_b[5071:5056];
  assign a_317 = io_a[5087:5072];
  assign b_317 = io_b[5087:5072];
  assign a_318 = io_a[5103:5088];
  assign b_318 = io_b[5103:5088];
  assign a_319 = io_a[5119:5104];
  assign b_319 = io_b[5119:5104];
  assign a_320 = io_a[5135:5120];
  assign b_320 = io_b[5135:5120];
  assign a_321 = io_a[5151:5136];
  assign b_321 = io_b[5151:5136];
  assign a_322 = io_a[5167:5152];
  assign b_322 = io_b[5167:5152];
  assign a_323 = io_a[5183:5168];
  assign b_323 = io_b[5183:5168];
  assign a_324 = io_a[5199:5184];
  assign b_324 = io_b[5199:5184];
  assign a_325 = io_a[5215:5200];
  assign b_325 = io_b[5215:5200];
  assign a_326 = io_a[5231:5216];
  assign b_326 = io_b[5231:5216];
  assign a_327 = io_a[5247:5232];
  assign b_327 = io_b[5247:5232];
  assign a_328 = io_a[5263:5248];
  assign b_328 = io_b[5263:5248];
  assign a_329 = io_a[5279:5264];
  assign b_329 = io_b[5279:5264];
  assign a_330 = io_a[5295:5280];
  assign b_330 = io_b[5295:5280];
  assign a_331 = io_a[5311:5296];
  assign b_331 = io_b[5311:5296];
  assign a_332 = io_a[5327:5312];
  assign b_332 = io_b[5327:5312];
  assign a_333 = io_a[5343:5328];
  assign b_333 = io_b[5343:5328];
  assign a_334 = io_a[5359:5344];
  assign b_334 = io_b[5359:5344];
  assign a_335 = io_a[5375:5360];
  assign b_335 = io_b[5375:5360];
  assign a_336 = io_a[5391:5376];
  assign b_336 = io_b[5391:5376];
  assign a_337 = io_a[5407:5392];
  assign b_337 = io_b[5407:5392];
  assign a_338 = io_a[5423:5408];
  assign b_338 = io_b[5423:5408];
  assign a_339 = io_a[5439:5424];
  assign b_339 = io_b[5439:5424];
  assign a_340 = io_a[5455:5440];
  assign b_340 = io_b[5455:5440];
  assign a_341 = io_a[5471:5456];
  assign b_341 = io_b[5471:5456];
  assign a_342 = io_a[5487:5472];
  assign b_342 = io_b[5487:5472];
  assign a_343 = io_a[5503:5488];
  assign b_343 = io_b[5503:5488];
  assign a_344 = io_a[5519:5504];
  assign b_344 = io_b[5519:5504];
  assign a_345 = io_a[5535:5520];
  assign b_345 = io_b[5535:5520];
  assign a_346 = io_a[5551:5536];
  assign b_346 = io_b[5551:5536];
  assign a_347 = io_a[5567:5552];
  assign b_347 = io_b[5567:5552];
  assign a_348 = io_a[5583:5568];
  assign b_348 = io_b[5583:5568];
  assign a_349 = io_a[5599:5584];
  assign b_349 = io_b[5599:5584];
  assign a_350 = io_a[5615:5600];
  assign b_350 = io_b[5615:5600];
  assign a_351 = io_a[5631:5616];
  assign b_351 = io_b[5631:5616];
  assign a_352 = io_a[5647:5632];
  assign b_352 = io_b[5647:5632];
  assign a_353 = io_a[5663:5648];
  assign b_353 = io_b[5663:5648];
  assign a_354 = io_a[5679:5664];
  assign b_354 = io_b[5679:5664];
  assign a_355 = io_a[5695:5680];
  assign b_355 = io_b[5695:5680];
  assign a_356 = io_a[5711:5696];
  assign b_356 = io_b[5711:5696];
  assign a_357 = io_a[5727:5712];
  assign b_357 = io_b[5727:5712];
  assign a_358 = io_a[5743:5728];
  assign b_358 = io_b[5743:5728];
  assign a_359 = io_a[5759:5744];
  assign b_359 = io_b[5759:5744];
  assign a_360 = io_a[5775:5760];
  assign b_360 = io_b[5775:5760];
  assign a_361 = io_a[5791:5776];
  assign b_361 = io_b[5791:5776];
  assign a_362 = io_a[5807:5792];
  assign b_362 = io_b[5807:5792];
  assign a_363 = io_a[5823:5808];
  assign b_363 = io_b[5823:5808];
  assign a_364 = io_a[5839:5824];
  assign b_364 = io_b[5839:5824];
  assign a_365 = io_a[5855:5840];
  assign b_365 = io_b[5855:5840];
  assign a_366 = io_a[5871:5856];
  assign b_366 = io_b[5871:5856];
  assign a_367 = io_a[5887:5872];
  assign b_367 = io_b[5887:5872];
  assign a_368 = io_a[5903:5888];
  assign b_368 = io_b[5903:5888];
  assign a_369 = io_a[5919:5904];
  assign b_369 = io_b[5919:5904];
  assign a_370 = io_a[5935:5920];
  assign b_370 = io_b[5935:5920];
  assign a_371 = io_a[5951:5936];
  assign b_371 = io_b[5951:5936];
  assign a_372 = io_a[5967:5952];
  assign b_372 = io_b[5967:5952];
  assign a_373 = io_a[5983:5968];
  assign b_373 = io_b[5983:5968];
  assign a_374 = io_a[5999:5984];
  assign b_374 = io_b[5999:5984];
  assign a_375 = io_a[6015:6000];
  assign b_375 = io_b[6015:6000];
  assign a_376 = io_a[6031:6016];
  assign b_376 = io_b[6031:6016];
  assign a_377 = io_a[6047:6032];
  assign b_377 = io_b[6047:6032];
  assign a_378 = io_a[6063:6048];
  assign b_378 = io_b[6063:6048];
  assign a_379 = io_a[6079:6064];
  assign b_379 = io_b[6079:6064];
  assign a_380 = io_a[6095:6080];
  assign b_380 = io_b[6095:6080];
  assign a_381 = io_a[6111:6096];
  assign b_381 = io_b[6111:6096];
  assign a_382 = io_a[6127:6112];
  assign b_382 = io_b[6127:6112];
  assign a_383 = io_a[6143:6128];
  assign b_383 = io_b[6143:6128];
  assign a_384 = io_a[6159:6144];
  assign b_384 = io_b[6159:6144];
  assign a_385 = io_a[6175:6160];
  assign b_385 = io_b[6175:6160];
  assign a_386 = io_a[6191:6176];
  assign b_386 = io_b[6191:6176];
  assign a_387 = io_a[6207:6192];
  assign b_387 = io_b[6207:6192];
  assign a_388 = io_a[6223:6208];
  assign b_388 = io_b[6223:6208];
  assign a_389 = io_a[6239:6224];
  assign b_389 = io_b[6239:6224];
  assign a_390 = io_a[6255:6240];
  assign b_390 = io_b[6255:6240];
  assign a_391 = io_a[6271:6256];
  assign b_391 = io_b[6271:6256];
  assign a_392 = io_a[6287:6272];
  assign b_392 = io_b[6287:6272];
  assign a_393 = io_a[6303:6288];
  assign b_393 = io_b[6303:6288];
  assign a_394 = io_a[6319:6304];
  assign b_394 = io_b[6319:6304];
  assign a_395 = io_a[6335:6320];
  assign b_395 = io_b[6335:6320];
  assign a_396 = io_a[6351:6336];
  assign b_396 = io_b[6351:6336];
  assign a_397 = io_a[6367:6352];
  assign b_397 = io_b[6367:6352];
  assign a_398 = io_a[6383:6368];
  assign b_398 = io_b[6383:6368];
  assign a_399 = io_a[6399:6384];
  assign b_399 = io_b[6399:6384];
  assign _T_803 = i == 9'h190;
  assign _T_804 = i != 9'h0;
  assign _GEN_1 = 9'h1 == i ? a_1 : a_0;
  assign _GEN_2 = 9'h2 == i ? a_2 : _GEN_1;
  assign _GEN_3 = 9'h3 == i ? a_3 : _GEN_2;
  assign _GEN_4 = 9'h4 == i ? a_4 : _GEN_3;
  assign _GEN_5 = 9'h5 == i ? a_5 : _GEN_4;
  assign _GEN_6 = 9'h6 == i ? a_6 : _GEN_5;
  assign _GEN_7 = 9'h7 == i ? a_7 : _GEN_6;
  assign _GEN_8 = 9'h8 == i ? a_8 : _GEN_7;
  assign _GEN_9 = 9'h9 == i ? a_9 : _GEN_8;
  assign _GEN_10 = 9'ha == i ? a_10 : _GEN_9;
  assign _GEN_11 = 9'hb == i ? a_11 : _GEN_10;
  assign _GEN_12 = 9'hc == i ? a_12 : _GEN_11;
  assign _GEN_13 = 9'hd == i ? a_13 : _GEN_12;
  assign _GEN_14 = 9'he == i ? a_14 : _GEN_13;
  assign _GEN_15 = 9'hf == i ? a_15 : _GEN_14;
  assign _GEN_16 = 9'h10 == i ? a_16 : _GEN_15;
  assign _GEN_17 = 9'h11 == i ? a_17 : _GEN_16;
  assign _GEN_18 = 9'h12 == i ? a_18 : _GEN_17;
  assign _GEN_19 = 9'h13 == i ? a_19 : _GEN_18;
  assign _GEN_20 = 9'h14 == i ? a_20 : _GEN_19;
  assign _GEN_21 = 9'h15 == i ? a_21 : _GEN_20;
  assign _GEN_22 = 9'h16 == i ? a_22 : _GEN_21;
  assign _GEN_23 = 9'h17 == i ? a_23 : _GEN_22;
  assign _GEN_24 = 9'h18 == i ? a_24 : _GEN_23;
  assign _GEN_25 = 9'h19 == i ? a_25 : _GEN_24;
  assign _GEN_26 = 9'h1a == i ? a_26 : _GEN_25;
  assign _GEN_27 = 9'h1b == i ? a_27 : _GEN_26;
  assign _GEN_28 = 9'h1c == i ? a_28 : _GEN_27;
  assign _GEN_29 = 9'h1d == i ? a_29 : _GEN_28;
  assign _GEN_30 = 9'h1e == i ? a_30 : _GEN_29;
  assign _GEN_31 = 9'h1f == i ? a_31 : _GEN_30;
  assign _GEN_32 = 9'h20 == i ? a_32 : _GEN_31;
  assign _GEN_33 = 9'h21 == i ? a_33 : _GEN_32;
  assign _GEN_34 = 9'h22 == i ? a_34 : _GEN_33;
  assign _GEN_35 = 9'h23 == i ? a_35 : _GEN_34;
  assign _GEN_36 = 9'h24 == i ? a_36 : _GEN_35;
  assign _GEN_37 = 9'h25 == i ? a_37 : _GEN_36;
  assign _GEN_38 = 9'h26 == i ? a_38 : _GEN_37;
  assign _GEN_39 = 9'h27 == i ? a_39 : _GEN_38;
  assign _GEN_40 = 9'h28 == i ? a_40 : _GEN_39;
  assign _GEN_41 = 9'h29 == i ? a_41 : _GEN_40;
  assign _GEN_42 = 9'h2a == i ? a_42 : _GEN_41;
  assign _GEN_43 = 9'h2b == i ? a_43 : _GEN_42;
  assign _GEN_44 = 9'h2c == i ? a_44 : _GEN_43;
  assign _GEN_45 = 9'h2d == i ? a_45 : _GEN_44;
  assign _GEN_46 = 9'h2e == i ? a_46 : _GEN_45;
  assign _GEN_47 = 9'h2f == i ? a_47 : _GEN_46;
  assign _GEN_48 = 9'h30 == i ? a_48 : _GEN_47;
  assign _GEN_49 = 9'h31 == i ? a_49 : _GEN_48;
  assign _GEN_50 = 9'h32 == i ? a_50 : _GEN_49;
  assign _GEN_51 = 9'h33 == i ? a_51 : _GEN_50;
  assign _GEN_52 = 9'h34 == i ? a_52 : _GEN_51;
  assign _GEN_53 = 9'h35 == i ? a_53 : _GEN_52;
  assign _GEN_54 = 9'h36 == i ? a_54 : _GEN_53;
  assign _GEN_55 = 9'h37 == i ? a_55 : _GEN_54;
  assign _GEN_56 = 9'h38 == i ? a_56 : _GEN_55;
  assign _GEN_57 = 9'h39 == i ? a_57 : _GEN_56;
  assign _GEN_58 = 9'h3a == i ? a_58 : _GEN_57;
  assign _GEN_59 = 9'h3b == i ? a_59 : _GEN_58;
  assign _GEN_60 = 9'h3c == i ? a_60 : _GEN_59;
  assign _GEN_61 = 9'h3d == i ? a_61 : _GEN_60;
  assign _GEN_62 = 9'h3e == i ? a_62 : _GEN_61;
  assign _GEN_63 = 9'h3f == i ? a_63 : _GEN_62;
  assign _GEN_64 = 9'h40 == i ? a_64 : _GEN_63;
  assign _GEN_65 = 9'h41 == i ? a_65 : _GEN_64;
  assign _GEN_66 = 9'h42 == i ? a_66 : _GEN_65;
  assign _GEN_67 = 9'h43 == i ? a_67 : _GEN_66;
  assign _GEN_68 = 9'h44 == i ? a_68 : _GEN_67;
  assign _GEN_69 = 9'h45 == i ? a_69 : _GEN_68;
  assign _GEN_70 = 9'h46 == i ? a_70 : _GEN_69;
  assign _GEN_71 = 9'h47 == i ? a_71 : _GEN_70;
  assign _GEN_72 = 9'h48 == i ? a_72 : _GEN_71;
  assign _GEN_73 = 9'h49 == i ? a_73 : _GEN_72;
  assign _GEN_74 = 9'h4a == i ? a_74 : _GEN_73;
  assign _GEN_75 = 9'h4b == i ? a_75 : _GEN_74;
  assign _GEN_76 = 9'h4c == i ? a_76 : _GEN_75;
  assign _GEN_77 = 9'h4d == i ? a_77 : _GEN_76;
  assign _GEN_78 = 9'h4e == i ? a_78 : _GEN_77;
  assign _GEN_79 = 9'h4f == i ? a_79 : _GEN_78;
  assign _GEN_80 = 9'h50 == i ? a_80 : _GEN_79;
  assign _GEN_81 = 9'h51 == i ? a_81 : _GEN_80;
  assign _GEN_82 = 9'h52 == i ? a_82 : _GEN_81;
  assign _GEN_83 = 9'h53 == i ? a_83 : _GEN_82;
  assign _GEN_84 = 9'h54 == i ? a_84 : _GEN_83;
  assign _GEN_85 = 9'h55 == i ? a_85 : _GEN_84;
  assign _GEN_86 = 9'h56 == i ? a_86 : _GEN_85;
  assign _GEN_87 = 9'h57 == i ? a_87 : _GEN_86;
  assign _GEN_88 = 9'h58 == i ? a_88 : _GEN_87;
  assign _GEN_89 = 9'h59 == i ? a_89 : _GEN_88;
  assign _GEN_90 = 9'h5a == i ? a_90 : _GEN_89;
  assign _GEN_91 = 9'h5b == i ? a_91 : _GEN_90;
  assign _GEN_92 = 9'h5c == i ? a_92 : _GEN_91;
  assign _GEN_93 = 9'h5d == i ? a_93 : _GEN_92;
  assign _GEN_94 = 9'h5e == i ? a_94 : _GEN_93;
  assign _GEN_95 = 9'h5f == i ? a_95 : _GEN_94;
  assign _GEN_96 = 9'h60 == i ? a_96 : _GEN_95;
  assign _GEN_97 = 9'h61 == i ? a_97 : _GEN_96;
  assign _GEN_98 = 9'h62 == i ? a_98 : _GEN_97;
  assign _GEN_99 = 9'h63 == i ? a_99 : _GEN_98;
  assign _GEN_100 = 9'h64 == i ? a_100 : _GEN_99;
  assign _GEN_101 = 9'h65 == i ? a_101 : _GEN_100;
  assign _GEN_102 = 9'h66 == i ? a_102 : _GEN_101;
  assign _GEN_103 = 9'h67 == i ? a_103 : _GEN_102;
  assign _GEN_104 = 9'h68 == i ? a_104 : _GEN_103;
  assign _GEN_105 = 9'h69 == i ? a_105 : _GEN_104;
  assign _GEN_106 = 9'h6a == i ? a_106 : _GEN_105;
  assign _GEN_107 = 9'h6b == i ? a_107 : _GEN_106;
  assign _GEN_108 = 9'h6c == i ? a_108 : _GEN_107;
  assign _GEN_109 = 9'h6d == i ? a_109 : _GEN_108;
  assign _GEN_110 = 9'h6e == i ? a_110 : _GEN_109;
  assign _GEN_111 = 9'h6f == i ? a_111 : _GEN_110;
  assign _GEN_112 = 9'h70 == i ? a_112 : _GEN_111;
  assign _GEN_113 = 9'h71 == i ? a_113 : _GEN_112;
  assign _GEN_114 = 9'h72 == i ? a_114 : _GEN_113;
  assign _GEN_115 = 9'h73 == i ? a_115 : _GEN_114;
  assign _GEN_116 = 9'h74 == i ? a_116 : _GEN_115;
  assign _GEN_117 = 9'h75 == i ? a_117 : _GEN_116;
  assign _GEN_118 = 9'h76 == i ? a_118 : _GEN_117;
  assign _GEN_119 = 9'h77 == i ? a_119 : _GEN_118;
  assign _GEN_120 = 9'h78 == i ? a_120 : _GEN_119;
  assign _GEN_121 = 9'h79 == i ? a_121 : _GEN_120;
  assign _GEN_122 = 9'h7a == i ? a_122 : _GEN_121;
  assign _GEN_123 = 9'h7b == i ? a_123 : _GEN_122;
  assign _GEN_124 = 9'h7c == i ? a_124 : _GEN_123;
  assign _GEN_125 = 9'h7d == i ? a_125 : _GEN_124;
  assign _GEN_126 = 9'h7e == i ? a_126 : _GEN_125;
  assign _GEN_127 = 9'h7f == i ? a_127 : _GEN_126;
  assign _GEN_128 = 9'h80 == i ? a_128 : _GEN_127;
  assign _GEN_129 = 9'h81 == i ? a_129 : _GEN_128;
  assign _GEN_130 = 9'h82 == i ? a_130 : _GEN_129;
  assign _GEN_131 = 9'h83 == i ? a_131 : _GEN_130;
  assign _GEN_132 = 9'h84 == i ? a_132 : _GEN_131;
  assign _GEN_133 = 9'h85 == i ? a_133 : _GEN_132;
  assign _GEN_134 = 9'h86 == i ? a_134 : _GEN_133;
  assign _GEN_135 = 9'h87 == i ? a_135 : _GEN_134;
  assign _GEN_136 = 9'h88 == i ? a_136 : _GEN_135;
  assign _GEN_137 = 9'h89 == i ? a_137 : _GEN_136;
  assign _GEN_138 = 9'h8a == i ? a_138 : _GEN_137;
  assign _GEN_139 = 9'h8b == i ? a_139 : _GEN_138;
  assign _GEN_140 = 9'h8c == i ? a_140 : _GEN_139;
  assign _GEN_141 = 9'h8d == i ? a_141 : _GEN_140;
  assign _GEN_142 = 9'h8e == i ? a_142 : _GEN_141;
  assign _GEN_143 = 9'h8f == i ? a_143 : _GEN_142;
  assign _GEN_144 = 9'h90 == i ? a_144 : _GEN_143;
  assign _GEN_145 = 9'h91 == i ? a_145 : _GEN_144;
  assign _GEN_146 = 9'h92 == i ? a_146 : _GEN_145;
  assign _GEN_147 = 9'h93 == i ? a_147 : _GEN_146;
  assign _GEN_148 = 9'h94 == i ? a_148 : _GEN_147;
  assign _GEN_149 = 9'h95 == i ? a_149 : _GEN_148;
  assign _GEN_150 = 9'h96 == i ? a_150 : _GEN_149;
  assign _GEN_151 = 9'h97 == i ? a_151 : _GEN_150;
  assign _GEN_152 = 9'h98 == i ? a_152 : _GEN_151;
  assign _GEN_153 = 9'h99 == i ? a_153 : _GEN_152;
  assign _GEN_154 = 9'h9a == i ? a_154 : _GEN_153;
  assign _GEN_155 = 9'h9b == i ? a_155 : _GEN_154;
  assign _GEN_156 = 9'h9c == i ? a_156 : _GEN_155;
  assign _GEN_157 = 9'h9d == i ? a_157 : _GEN_156;
  assign _GEN_158 = 9'h9e == i ? a_158 : _GEN_157;
  assign _GEN_159 = 9'h9f == i ? a_159 : _GEN_158;
  assign _GEN_160 = 9'ha0 == i ? a_160 : _GEN_159;
  assign _GEN_161 = 9'ha1 == i ? a_161 : _GEN_160;
  assign _GEN_162 = 9'ha2 == i ? a_162 : _GEN_161;
  assign _GEN_163 = 9'ha3 == i ? a_163 : _GEN_162;
  assign _GEN_164 = 9'ha4 == i ? a_164 : _GEN_163;
  assign _GEN_165 = 9'ha5 == i ? a_165 : _GEN_164;
  assign _GEN_166 = 9'ha6 == i ? a_166 : _GEN_165;
  assign _GEN_167 = 9'ha7 == i ? a_167 : _GEN_166;
  assign _GEN_168 = 9'ha8 == i ? a_168 : _GEN_167;
  assign _GEN_169 = 9'ha9 == i ? a_169 : _GEN_168;
  assign _GEN_170 = 9'haa == i ? a_170 : _GEN_169;
  assign _GEN_171 = 9'hab == i ? a_171 : _GEN_170;
  assign _GEN_172 = 9'hac == i ? a_172 : _GEN_171;
  assign _GEN_173 = 9'had == i ? a_173 : _GEN_172;
  assign _GEN_174 = 9'hae == i ? a_174 : _GEN_173;
  assign _GEN_175 = 9'haf == i ? a_175 : _GEN_174;
  assign _GEN_176 = 9'hb0 == i ? a_176 : _GEN_175;
  assign _GEN_177 = 9'hb1 == i ? a_177 : _GEN_176;
  assign _GEN_178 = 9'hb2 == i ? a_178 : _GEN_177;
  assign _GEN_179 = 9'hb3 == i ? a_179 : _GEN_178;
  assign _GEN_180 = 9'hb4 == i ? a_180 : _GEN_179;
  assign _GEN_181 = 9'hb5 == i ? a_181 : _GEN_180;
  assign _GEN_182 = 9'hb6 == i ? a_182 : _GEN_181;
  assign _GEN_183 = 9'hb7 == i ? a_183 : _GEN_182;
  assign _GEN_184 = 9'hb8 == i ? a_184 : _GEN_183;
  assign _GEN_185 = 9'hb9 == i ? a_185 : _GEN_184;
  assign _GEN_186 = 9'hba == i ? a_186 : _GEN_185;
  assign _GEN_187 = 9'hbb == i ? a_187 : _GEN_186;
  assign _GEN_188 = 9'hbc == i ? a_188 : _GEN_187;
  assign _GEN_189 = 9'hbd == i ? a_189 : _GEN_188;
  assign _GEN_190 = 9'hbe == i ? a_190 : _GEN_189;
  assign _GEN_191 = 9'hbf == i ? a_191 : _GEN_190;
  assign _GEN_192 = 9'hc0 == i ? a_192 : _GEN_191;
  assign _GEN_193 = 9'hc1 == i ? a_193 : _GEN_192;
  assign _GEN_194 = 9'hc2 == i ? a_194 : _GEN_193;
  assign _GEN_195 = 9'hc3 == i ? a_195 : _GEN_194;
  assign _GEN_196 = 9'hc4 == i ? a_196 : _GEN_195;
  assign _GEN_197 = 9'hc5 == i ? a_197 : _GEN_196;
  assign _GEN_198 = 9'hc6 == i ? a_198 : _GEN_197;
  assign _GEN_199 = 9'hc7 == i ? a_199 : _GEN_198;
  assign _GEN_200 = 9'hc8 == i ? a_200 : _GEN_199;
  assign _GEN_201 = 9'hc9 == i ? a_201 : _GEN_200;
  assign _GEN_202 = 9'hca == i ? a_202 : _GEN_201;
  assign _GEN_203 = 9'hcb == i ? a_203 : _GEN_202;
  assign _GEN_204 = 9'hcc == i ? a_204 : _GEN_203;
  assign _GEN_205 = 9'hcd == i ? a_205 : _GEN_204;
  assign _GEN_206 = 9'hce == i ? a_206 : _GEN_205;
  assign _GEN_207 = 9'hcf == i ? a_207 : _GEN_206;
  assign _GEN_208 = 9'hd0 == i ? a_208 : _GEN_207;
  assign _GEN_209 = 9'hd1 == i ? a_209 : _GEN_208;
  assign _GEN_210 = 9'hd2 == i ? a_210 : _GEN_209;
  assign _GEN_211 = 9'hd3 == i ? a_211 : _GEN_210;
  assign _GEN_212 = 9'hd4 == i ? a_212 : _GEN_211;
  assign _GEN_213 = 9'hd5 == i ? a_213 : _GEN_212;
  assign _GEN_214 = 9'hd6 == i ? a_214 : _GEN_213;
  assign _GEN_215 = 9'hd7 == i ? a_215 : _GEN_214;
  assign _GEN_216 = 9'hd8 == i ? a_216 : _GEN_215;
  assign _GEN_217 = 9'hd9 == i ? a_217 : _GEN_216;
  assign _GEN_218 = 9'hda == i ? a_218 : _GEN_217;
  assign _GEN_219 = 9'hdb == i ? a_219 : _GEN_218;
  assign _GEN_220 = 9'hdc == i ? a_220 : _GEN_219;
  assign _GEN_221 = 9'hdd == i ? a_221 : _GEN_220;
  assign _GEN_222 = 9'hde == i ? a_222 : _GEN_221;
  assign _GEN_223 = 9'hdf == i ? a_223 : _GEN_222;
  assign _GEN_224 = 9'he0 == i ? a_224 : _GEN_223;
  assign _GEN_225 = 9'he1 == i ? a_225 : _GEN_224;
  assign _GEN_226 = 9'he2 == i ? a_226 : _GEN_225;
  assign _GEN_227 = 9'he3 == i ? a_227 : _GEN_226;
  assign _GEN_228 = 9'he4 == i ? a_228 : _GEN_227;
  assign _GEN_229 = 9'he5 == i ? a_229 : _GEN_228;
  assign _GEN_230 = 9'he6 == i ? a_230 : _GEN_229;
  assign _GEN_231 = 9'he7 == i ? a_231 : _GEN_230;
  assign _GEN_232 = 9'he8 == i ? a_232 : _GEN_231;
  assign _GEN_233 = 9'he9 == i ? a_233 : _GEN_232;
  assign _GEN_234 = 9'hea == i ? a_234 : _GEN_233;
  assign _GEN_235 = 9'heb == i ? a_235 : _GEN_234;
  assign _GEN_236 = 9'hec == i ? a_236 : _GEN_235;
  assign _GEN_237 = 9'hed == i ? a_237 : _GEN_236;
  assign _GEN_238 = 9'hee == i ? a_238 : _GEN_237;
  assign _GEN_239 = 9'hef == i ? a_239 : _GEN_238;
  assign _GEN_240 = 9'hf0 == i ? a_240 : _GEN_239;
  assign _GEN_241 = 9'hf1 == i ? a_241 : _GEN_240;
  assign _GEN_242 = 9'hf2 == i ? a_242 : _GEN_241;
  assign _GEN_243 = 9'hf3 == i ? a_243 : _GEN_242;
  assign _GEN_244 = 9'hf4 == i ? a_244 : _GEN_243;
  assign _GEN_245 = 9'hf5 == i ? a_245 : _GEN_244;
  assign _GEN_246 = 9'hf6 == i ? a_246 : _GEN_245;
  assign _GEN_247 = 9'hf7 == i ? a_247 : _GEN_246;
  assign _GEN_248 = 9'hf8 == i ? a_248 : _GEN_247;
  assign _GEN_249 = 9'hf9 == i ? a_249 : _GEN_248;
  assign _GEN_250 = 9'hfa == i ? a_250 : _GEN_249;
  assign _GEN_251 = 9'hfb == i ? a_251 : _GEN_250;
  assign _GEN_252 = 9'hfc == i ? a_252 : _GEN_251;
  assign _GEN_253 = 9'hfd == i ? a_253 : _GEN_252;
  assign _GEN_254 = 9'hfe == i ? a_254 : _GEN_253;
  assign _GEN_255 = 9'hff == i ? a_255 : _GEN_254;
  assign _GEN_256 = 9'h100 == i ? a_256 : _GEN_255;
  assign _GEN_257 = 9'h101 == i ? a_257 : _GEN_256;
  assign _GEN_258 = 9'h102 == i ? a_258 : _GEN_257;
  assign _GEN_259 = 9'h103 == i ? a_259 : _GEN_258;
  assign _GEN_260 = 9'h104 == i ? a_260 : _GEN_259;
  assign _GEN_261 = 9'h105 == i ? a_261 : _GEN_260;
  assign _GEN_262 = 9'h106 == i ? a_262 : _GEN_261;
  assign _GEN_263 = 9'h107 == i ? a_263 : _GEN_262;
  assign _GEN_264 = 9'h108 == i ? a_264 : _GEN_263;
  assign _GEN_265 = 9'h109 == i ? a_265 : _GEN_264;
  assign _GEN_266 = 9'h10a == i ? a_266 : _GEN_265;
  assign _GEN_267 = 9'h10b == i ? a_267 : _GEN_266;
  assign _GEN_268 = 9'h10c == i ? a_268 : _GEN_267;
  assign _GEN_269 = 9'h10d == i ? a_269 : _GEN_268;
  assign _GEN_270 = 9'h10e == i ? a_270 : _GEN_269;
  assign _GEN_271 = 9'h10f == i ? a_271 : _GEN_270;
  assign _GEN_272 = 9'h110 == i ? a_272 : _GEN_271;
  assign _GEN_273 = 9'h111 == i ? a_273 : _GEN_272;
  assign _GEN_274 = 9'h112 == i ? a_274 : _GEN_273;
  assign _GEN_275 = 9'h113 == i ? a_275 : _GEN_274;
  assign _GEN_276 = 9'h114 == i ? a_276 : _GEN_275;
  assign _GEN_277 = 9'h115 == i ? a_277 : _GEN_276;
  assign _GEN_278 = 9'h116 == i ? a_278 : _GEN_277;
  assign _GEN_279 = 9'h117 == i ? a_279 : _GEN_278;
  assign _GEN_280 = 9'h118 == i ? a_280 : _GEN_279;
  assign _GEN_281 = 9'h119 == i ? a_281 : _GEN_280;
  assign _GEN_282 = 9'h11a == i ? a_282 : _GEN_281;
  assign _GEN_283 = 9'h11b == i ? a_283 : _GEN_282;
  assign _GEN_284 = 9'h11c == i ? a_284 : _GEN_283;
  assign _GEN_285 = 9'h11d == i ? a_285 : _GEN_284;
  assign _GEN_286 = 9'h11e == i ? a_286 : _GEN_285;
  assign _GEN_287 = 9'h11f == i ? a_287 : _GEN_286;
  assign _GEN_288 = 9'h120 == i ? a_288 : _GEN_287;
  assign _GEN_289 = 9'h121 == i ? a_289 : _GEN_288;
  assign _GEN_290 = 9'h122 == i ? a_290 : _GEN_289;
  assign _GEN_291 = 9'h123 == i ? a_291 : _GEN_290;
  assign _GEN_292 = 9'h124 == i ? a_292 : _GEN_291;
  assign _GEN_293 = 9'h125 == i ? a_293 : _GEN_292;
  assign _GEN_294 = 9'h126 == i ? a_294 : _GEN_293;
  assign _GEN_295 = 9'h127 == i ? a_295 : _GEN_294;
  assign _GEN_296 = 9'h128 == i ? a_296 : _GEN_295;
  assign _GEN_297 = 9'h129 == i ? a_297 : _GEN_296;
  assign _GEN_298 = 9'h12a == i ? a_298 : _GEN_297;
  assign _GEN_299 = 9'h12b == i ? a_299 : _GEN_298;
  assign _GEN_300 = 9'h12c == i ? a_300 : _GEN_299;
  assign _GEN_301 = 9'h12d == i ? a_301 : _GEN_300;
  assign _GEN_302 = 9'h12e == i ? a_302 : _GEN_301;
  assign _GEN_303 = 9'h12f == i ? a_303 : _GEN_302;
  assign _GEN_304 = 9'h130 == i ? a_304 : _GEN_303;
  assign _GEN_305 = 9'h131 == i ? a_305 : _GEN_304;
  assign _GEN_306 = 9'h132 == i ? a_306 : _GEN_305;
  assign _GEN_307 = 9'h133 == i ? a_307 : _GEN_306;
  assign _GEN_308 = 9'h134 == i ? a_308 : _GEN_307;
  assign _GEN_309 = 9'h135 == i ? a_309 : _GEN_308;
  assign _GEN_310 = 9'h136 == i ? a_310 : _GEN_309;
  assign _GEN_311 = 9'h137 == i ? a_311 : _GEN_310;
  assign _GEN_312 = 9'h138 == i ? a_312 : _GEN_311;
  assign _GEN_313 = 9'h139 == i ? a_313 : _GEN_312;
  assign _GEN_314 = 9'h13a == i ? a_314 : _GEN_313;
  assign _GEN_315 = 9'h13b == i ? a_315 : _GEN_314;
  assign _GEN_316 = 9'h13c == i ? a_316 : _GEN_315;
  assign _GEN_317 = 9'h13d == i ? a_317 : _GEN_316;
  assign _GEN_318 = 9'h13e == i ? a_318 : _GEN_317;
  assign _GEN_319 = 9'h13f == i ? a_319 : _GEN_318;
  assign _GEN_320 = 9'h140 == i ? a_320 : _GEN_319;
  assign _GEN_321 = 9'h141 == i ? a_321 : _GEN_320;
  assign _GEN_322 = 9'h142 == i ? a_322 : _GEN_321;
  assign _GEN_323 = 9'h143 == i ? a_323 : _GEN_322;
  assign _GEN_324 = 9'h144 == i ? a_324 : _GEN_323;
  assign _GEN_325 = 9'h145 == i ? a_325 : _GEN_324;
  assign _GEN_326 = 9'h146 == i ? a_326 : _GEN_325;
  assign _GEN_327 = 9'h147 == i ? a_327 : _GEN_326;
  assign _GEN_328 = 9'h148 == i ? a_328 : _GEN_327;
  assign _GEN_329 = 9'h149 == i ? a_329 : _GEN_328;
  assign _GEN_330 = 9'h14a == i ? a_330 : _GEN_329;
  assign _GEN_331 = 9'h14b == i ? a_331 : _GEN_330;
  assign _GEN_332 = 9'h14c == i ? a_332 : _GEN_331;
  assign _GEN_333 = 9'h14d == i ? a_333 : _GEN_332;
  assign _GEN_334 = 9'h14e == i ? a_334 : _GEN_333;
  assign _GEN_335 = 9'h14f == i ? a_335 : _GEN_334;
  assign _GEN_336 = 9'h150 == i ? a_336 : _GEN_335;
  assign _GEN_337 = 9'h151 == i ? a_337 : _GEN_336;
  assign _GEN_338 = 9'h152 == i ? a_338 : _GEN_337;
  assign _GEN_339 = 9'h153 == i ? a_339 : _GEN_338;
  assign _GEN_340 = 9'h154 == i ? a_340 : _GEN_339;
  assign _GEN_341 = 9'h155 == i ? a_341 : _GEN_340;
  assign _GEN_342 = 9'h156 == i ? a_342 : _GEN_341;
  assign _GEN_343 = 9'h157 == i ? a_343 : _GEN_342;
  assign _GEN_344 = 9'h158 == i ? a_344 : _GEN_343;
  assign _GEN_345 = 9'h159 == i ? a_345 : _GEN_344;
  assign _GEN_346 = 9'h15a == i ? a_346 : _GEN_345;
  assign _GEN_347 = 9'h15b == i ? a_347 : _GEN_346;
  assign _GEN_348 = 9'h15c == i ? a_348 : _GEN_347;
  assign _GEN_349 = 9'h15d == i ? a_349 : _GEN_348;
  assign _GEN_350 = 9'h15e == i ? a_350 : _GEN_349;
  assign _GEN_351 = 9'h15f == i ? a_351 : _GEN_350;
  assign _GEN_352 = 9'h160 == i ? a_352 : _GEN_351;
  assign _GEN_353 = 9'h161 == i ? a_353 : _GEN_352;
  assign _GEN_354 = 9'h162 == i ? a_354 : _GEN_353;
  assign _GEN_355 = 9'h163 == i ? a_355 : _GEN_354;
  assign _GEN_356 = 9'h164 == i ? a_356 : _GEN_355;
  assign _GEN_357 = 9'h165 == i ? a_357 : _GEN_356;
  assign _GEN_358 = 9'h166 == i ? a_358 : _GEN_357;
  assign _GEN_359 = 9'h167 == i ? a_359 : _GEN_358;
  assign _GEN_360 = 9'h168 == i ? a_360 : _GEN_359;
  assign _GEN_361 = 9'h169 == i ? a_361 : _GEN_360;
  assign _GEN_362 = 9'h16a == i ? a_362 : _GEN_361;
  assign _GEN_363 = 9'h16b == i ? a_363 : _GEN_362;
  assign _GEN_364 = 9'h16c == i ? a_364 : _GEN_363;
  assign _GEN_365 = 9'h16d == i ? a_365 : _GEN_364;
  assign _GEN_366 = 9'h16e == i ? a_366 : _GEN_365;
  assign _GEN_367 = 9'h16f == i ? a_367 : _GEN_366;
  assign _GEN_368 = 9'h170 == i ? a_368 : _GEN_367;
  assign _GEN_369 = 9'h171 == i ? a_369 : _GEN_368;
  assign _GEN_370 = 9'h172 == i ? a_370 : _GEN_369;
  assign _GEN_371 = 9'h173 == i ? a_371 : _GEN_370;
  assign _GEN_372 = 9'h174 == i ? a_372 : _GEN_371;
  assign _GEN_373 = 9'h175 == i ? a_373 : _GEN_372;
  assign _GEN_374 = 9'h176 == i ? a_374 : _GEN_373;
  assign _GEN_375 = 9'h177 == i ? a_375 : _GEN_374;
  assign _GEN_376 = 9'h178 == i ? a_376 : _GEN_375;
  assign _GEN_377 = 9'h179 == i ? a_377 : _GEN_376;
  assign _GEN_378 = 9'h17a == i ? a_378 : _GEN_377;
  assign _GEN_379 = 9'h17b == i ? a_379 : _GEN_378;
  assign _GEN_380 = 9'h17c == i ? a_380 : _GEN_379;
  assign _GEN_381 = 9'h17d == i ? a_381 : _GEN_380;
  assign _GEN_382 = 9'h17e == i ? a_382 : _GEN_381;
  assign _GEN_383 = 9'h17f == i ? a_383 : _GEN_382;
  assign _GEN_384 = 9'h180 == i ? a_384 : _GEN_383;
  assign _GEN_385 = 9'h181 == i ? a_385 : _GEN_384;
  assign _GEN_386 = 9'h182 == i ? a_386 : _GEN_385;
  assign _GEN_387 = 9'h183 == i ? a_387 : _GEN_386;
  assign _GEN_388 = 9'h184 == i ? a_388 : _GEN_387;
  assign _GEN_389 = 9'h185 == i ? a_389 : _GEN_388;
  assign _GEN_390 = 9'h186 == i ? a_390 : _GEN_389;
  assign _GEN_391 = 9'h187 == i ? a_391 : _GEN_390;
  assign _GEN_392 = 9'h188 == i ? a_392 : _GEN_391;
  assign _GEN_393 = 9'h189 == i ? a_393 : _GEN_392;
  assign _GEN_394 = 9'h18a == i ? a_394 : _GEN_393;
  assign _GEN_395 = 9'h18b == i ? a_395 : _GEN_394;
  assign _GEN_396 = 9'h18c == i ? a_396 : _GEN_395;
  assign _GEN_397 = 9'h18d == i ? a_397 : _GEN_396;
  assign _GEN_398 = 9'h18e == i ? a_398 : _GEN_397;
  assign _GEN_399 = 9'h18f == i ? a_399 : _GEN_398;
  assign _GEN_401 = 9'h1 == i ? b_1 : b_0;
  assign _GEN_402 = 9'h2 == i ? b_2 : _GEN_401;
  assign _GEN_403 = 9'h3 == i ? b_3 : _GEN_402;
  assign _GEN_404 = 9'h4 == i ? b_4 : _GEN_403;
  assign _GEN_405 = 9'h5 == i ? b_5 : _GEN_404;
  assign _GEN_406 = 9'h6 == i ? b_6 : _GEN_405;
  assign _GEN_407 = 9'h7 == i ? b_7 : _GEN_406;
  assign _GEN_408 = 9'h8 == i ? b_8 : _GEN_407;
  assign _GEN_409 = 9'h9 == i ? b_9 : _GEN_408;
  assign _GEN_410 = 9'ha == i ? b_10 : _GEN_409;
  assign _GEN_411 = 9'hb == i ? b_11 : _GEN_410;
  assign _GEN_412 = 9'hc == i ? b_12 : _GEN_411;
  assign _GEN_413 = 9'hd == i ? b_13 : _GEN_412;
  assign _GEN_414 = 9'he == i ? b_14 : _GEN_413;
  assign _GEN_415 = 9'hf == i ? b_15 : _GEN_414;
  assign _GEN_416 = 9'h10 == i ? b_16 : _GEN_415;
  assign _GEN_417 = 9'h11 == i ? b_17 : _GEN_416;
  assign _GEN_418 = 9'h12 == i ? b_18 : _GEN_417;
  assign _GEN_419 = 9'h13 == i ? b_19 : _GEN_418;
  assign _GEN_420 = 9'h14 == i ? b_20 : _GEN_419;
  assign _GEN_421 = 9'h15 == i ? b_21 : _GEN_420;
  assign _GEN_422 = 9'h16 == i ? b_22 : _GEN_421;
  assign _GEN_423 = 9'h17 == i ? b_23 : _GEN_422;
  assign _GEN_424 = 9'h18 == i ? b_24 : _GEN_423;
  assign _GEN_425 = 9'h19 == i ? b_25 : _GEN_424;
  assign _GEN_426 = 9'h1a == i ? b_26 : _GEN_425;
  assign _GEN_427 = 9'h1b == i ? b_27 : _GEN_426;
  assign _GEN_428 = 9'h1c == i ? b_28 : _GEN_427;
  assign _GEN_429 = 9'h1d == i ? b_29 : _GEN_428;
  assign _GEN_430 = 9'h1e == i ? b_30 : _GEN_429;
  assign _GEN_431 = 9'h1f == i ? b_31 : _GEN_430;
  assign _GEN_432 = 9'h20 == i ? b_32 : _GEN_431;
  assign _GEN_433 = 9'h21 == i ? b_33 : _GEN_432;
  assign _GEN_434 = 9'h22 == i ? b_34 : _GEN_433;
  assign _GEN_435 = 9'h23 == i ? b_35 : _GEN_434;
  assign _GEN_436 = 9'h24 == i ? b_36 : _GEN_435;
  assign _GEN_437 = 9'h25 == i ? b_37 : _GEN_436;
  assign _GEN_438 = 9'h26 == i ? b_38 : _GEN_437;
  assign _GEN_439 = 9'h27 == i ? b_39 : _GEN_438;
  assign _GEN_440 = 9'h28 == i ? b_40 : _GEN_439;
  assign _GEN_441 = 9'h29 == i ? b_41 : _GEN_440;
  assign _GEN_442 = 9'h2a == i ? b_42 : _GEN_441;
  assign _GEN_443 = 9'h2b == i ? b_43 : _GEN_442;
  assign _GEN_444 = 9'h2c == i ? b_44 : _GEN_443;
  assign _GEN_445 = 9'h2d == i ? b_45 : _GEN_444;
  assign _GEN_446 = 9'h2e == i ? b_46 : _GEN_445;
  assign _GEN_447 = 9'h2f == i ? b_47 : _GEN_446;
  assign _GEN_448 = 9'h30 == i ? b_48 : _GEN_447;
  assign _GEN_449 = 9'h31 == i ? b_49 : _GEN_448;
  assign _GEN_450 = 9'h32 == i ? b_50 : _GEN_449;
  assign _GEN_451 = 9'h33 == i ? b_51 : _GEN_450;
  assign _GEN_452 = 9'h34 == i ? b_52 : _GEN_451;
  assign _GEN_453 = 9'h35 == i ? b_53 : _GEN_452;
  assign _GEN_454 = 9'h36 == i ? b_54 : _GEN_453;
  assign _GEN_455 = 9'h37 == i ? b_55 : _GEN_454;
  assign _GEN_456 = 9'h38 == i ? b_56 : _GEN_455;
  assign _GEN_457 = 9'h39 == i ? b_57 : _GEN_456;
  assign _GEN_458 = 9'h3a == i ? b_58 : _GEN_457;
  assign _GEN_459 = 9'h3b == i ? b_59 : _GEN_458;
  assign _GEN_460 = 9'h3c == i ? b_60 : _GEN_459;
  assign _GEN_461 = 9'h3d == i ? b_61 : _GEN_460;
  assign _GEN_462 = 9'h3e == i ? b_62 : _GEN_461;
  assign _GEN_463 = 9'h3f == i ? b_63 : _GEN_462;
  assign _GEN_464 = 9'h40 == i ? b_64 : _GEN_463;
  assign _GEN_465 = 9'h41 == i ? b_65 : _GEN_464;
  assign _GEN_466 = 9'h42 == i ? b_66 : _GEN_465;
  assign _GEN_467 = 9'h43 == i ? b_67 : _GEN_466;
  assign _GEN_468 = 9'h44 == i ? b_68 : _GEN_467;
  assign _GEN_469 = 9'h45 == i ? b_69 : _GEN_468;
  assign _GEN_470 = 9'h46 == i ? b_70 : _GEN_469;
  assign _GEN_471 = 9'h47 == i ? b_71 : _GEN_470;
  assign _GEN_472 = 9'h48 == i ? b_72 : _GEN_471;
  assign _GEN_473 = 9'h49 == i ? b_73 : _GEN_472;
  assign _GEN_474 = 9'h4a == i ? b_74 : _GEN_473;
  assign _GEN_475 = 9'h4b == i ? b_75 : _GEN_474;
  assign _GEN_476 = 9'h4c == i ? b_76 : _GEN_475;
  assign _GEN_477 = 9'h4d == i ? b_77 : _GEN_476;
  assign _GEN_478 = 9'h4e == i ? b_78 : _GEN_477;
  assign _GEN_479 = 9'h4f == i ? b_79 : _GEN_478;
  assign _GEN_480 = 9'h50 == i ? b_80 : _GEN_479;
  assign _GEN_481 = 9'h51 == i ? b_81 : _GEN_480;
  assign _GEN_482 = 9'h52 == i ? b_82 : _GEN_481;
  assign _GEN_483 = 9'h53 == i ? b_83 : _GEN_482;
  assign _GEN_484 = 9'h54 == i ? b_84 : _GEN_483;
  assign _GEN_485 = 9'h55 == i ? b_85 : _GEN_484;
  assign _GEN_486 = 9'h56 == i ? b_86 : _GEN_485;
  assign _GEN_487 = 9'h57 == i ? b_87 : _GEN_486;
  assign _GEN_488 = 9'h58 == i ? b_88 : _GEN_487;
  assign _GEN_489 = 9'h59 == i ? b_89 : _GEN_488;
  assign _GEN_490 = 9'h5a == i ? b_90 : _GEN_489;
  assign _GEN_491 = 9'h5b == i ? b_91 : _GEN_490;
  assign _GEN_492 = 9'h5c == i ? b_92 : _GEN_491;
  assign _GEN_493 = 9'h5d == i ? b_93 : _GEN_492;
  assign _GEN_494 = 9'h5e == i ? b_94 : _GEN_493;
  assign _GEN_495 = 9'h5f == i ? b_95 : _GEN_494;
  assign _GEN_496 = 9'h60 == i ? b_96 : _GEN_495;
  assign _GEN_497 = 9'h61 == i ? b_97 : _GEN_496;
  assign _GEN_498 = 9'h62 == i ? b_98 : _GEN_497;
  assign _GEN_499 = 9'h63 == i ? b_99 : _GEN_498;
  assign _GEN_500 = 9'h64 == i ? b_100 : _GEN_499;
  assign _GEN_501 = 9'h65 == i ? b_101 : _GEN_500;
  assign _GEN_502 = 9'h66 == i ? b_102 : _GEN_501;
  assign _GEN_503 = 9'h67 == i ? b_103 : _GEN_502;
  assign _GEN_504 = 9'h68 == i ? b_104 : _GEN_503;
  assign _GEN_505 = 9'h69 == i ? b_105 : _GEN_504;
  assign _GEN_506 = 9'h6a == i ? b_106 : _GEN_505;
  assign _GEN_507 = 9'h6b == i ? b_107 : _GEN_506;
  assign _GEN_508 = 9'h6c == i ? b_108 : _GEN_507;
  assign _GEN_509 = 9'h6d == i ? b_109 : _GEN_508;
  assign _GEN_510 = 9'h6e == i ? b_110 : _GEN_509;
  assign _GEN_511 = 9'h6f == i ? b_111 : _GEN_510;
  assign _GEN_512 = 9'h70 == i ? b_112 : _GEN_511;
  assign _GEN_513 = 9'h71 == i ? b_113 : _GEN_512;
  assign _GEN_514 = 9'h72 == i ? b_114 : _GEN_513;
  assign _GEN_515 = 9'h73 == i ? b_115 : _GEN_514;
  assign _GEN_516 = 9'h74 == i ? b_116 : _GEN_515;
  assign _GEN_517 = 9'h75 == i ? b_117 : _GEN_516;
  assign _GEN_518 = 9'h76 == i ? b_118 : _GEN_517;
  assign _GEN_519 = 9'h77 == i ? b_119 : _GEN_518;
  assign _GEN_520 = 9'h78 == i ? b_120 : _GEN_519;
  assign _GEN_521 = 9'h79 == i ? b_121 : _GEN_520;
  assign _GEN_522 = 9'h7a == i ? b_122 : _GEN_521;
  assign _GEN_523 = 9'h7b == i ? b_123 : _GEN_522;
  assign _GEN_524 = 9'h7c == i ? b_124 : _GEN_523;
  assign _GEN_525 = 9'h7d == i ? b_125 : _GEN_524;
  assign _GEN_526 = 9'h7e == i ? b_126 : _GEN_525;
  assign _GEN_527 = 9'h7f == i ? b_127 : _GEN_526;
  assign _GEN_528 = 9'h80 == i ? b_128 : _GEN_527;
  assign _GEN_529 = 9'h81 == i ? b_129 : _GEN_528;
  assign _GEN_530 = 9'h82 == i ? b_130 : _GEN_529;
  assign _GEN_531 = 9'h83 == i ? b_131 : _GEN_530;
  assign _GEN_532 = 9'h84 == i ? b_132 : _GEN_531;
  assign _GEN_533 = 9'h85 == i ? b_133 : _GEN_532;
  assign _GEN_534 = 9'h86 == i ? b_134 : _GEN_533;
  assign _GEN_535 = 9'h87 == i ? b_135 : _GEN_534;
  assign _GEN_536 = 9'h88 == i ? b_136 : _GEN_535;
  assign _GEN_537 = 9'h89 == i ? b_137 : _GEN_536;
  assign _GEN_538 = 9'h8a == i ? b_138 : _GEN_537;
  assign _GEN_539 = 9'h8b == i ? b_139 : _GEN_538;
  assign _GEN_540 = 9'h8c == i ? b_140 : _GEN_539;
  assign _GEN_541 = 9'h8d == i ? b_141 : _GEN_540;
  assign _GEN_542 = 9'h8e == i ? b_142 : _GEN_541;
  assign _GEN_543 = 9'h8f == i ? b_143 : _GEN_542;
  assign _GEN_544 = 9'h90 == i ? b_144 : _GEN_543;
  assign _GEN_545 = 9'h91 == i ? b_145 : _GEN_544;
  assign _GEN_546 = 9'h92 == i ? b_146 : _GEN_545;
  assign _GEN_547 = 9'h93 == i ? b_147 : _GEN_546;
  assign _GEN_548 = 9'h94 == i ? b_148 : _GEN_547;
  assign _GEN_549 = 9'h95 == i ? b_149 : _GEN_548;
  assign _GEN_550 = 9'h96 == i ? b_150 : _GEN_549;
  assign _GEN_551 = 9'h97 == i ? b_151 : _GEN_550;
  assign _GEN_552 = 9'h98 == i ? b_152 : _GEN_551;
  assign _GEN_553 = 9'h99 == i ? b_153 : _GEN_552;
  assign _GEN_554 = 9'h9a == i ? b_154 : _GEN_553;
  assign _GEN_555 = 9'h9b == i ? b_155 : _GEN_554;
  assign _GEN_556 = 9'h9c == i ? b_156 : _GEN_555;
  assign _GEN_557 = 9'h9d == i ? b_157 : _GEN_556;
  assign _GEN_558 = 9'h9e == i ? b_158 : _GEN_557;
  assign _GEN_559 = 9'h9f == i ? b_159 : _GEN_558;
  assign _GEN_560 = 9'ha0 == i ? b_160 : _GEN_559;
  assign _GEN_561 = 9'ha1 == i ? b_161 : _GEN_560;
  assign _GEN_562 = 9'ha2 == i ? b_162 : _GEN_561;
  assign _GEN_563 = 9'ha3 == i ? b_163 : _GEN_562;
  assign _GEN_564 = 9'ha4 == i ? b_164 : _GEN_563;
  assign _GEN_565 = 9'ha5 == i ? b_165 : _GEN_564;
  assign _GEN_566 = 9'ha6 == i ? b_166 : _GEN_565;
  assign _GEN_567 = 9'ha7 == i ? b_167 : _GEN_566;
  assign _GEN_568 = 9'ha8 == i ? b_168 : _GEN_567;
  assign _GEN_569 = 9'ha9 == i ? b_169 : _GEN_568;
  assign _GEN_570 = 9'haa == i ? b_170 : _GEN_569;
  assign _GEN_571 = 9'hab == i ? b_171 : _GEN_570;
  assign _GEN_572 = 9'hac == i ? b_172 : _GEN_571;
  assign _GEN_573 = 9'had == i ? b_173 : _GEN_572;
  assign _GEN_574 = 9'hae == i ? b_174 : _GEN_573;
  assign _GEN_575 = 9'haf == i ? b_175 : _GEN_574;
  assign _GEN_576 = 9'hb0 == i ? b_176 : _GEN_575;
  assign _GEN_577 = 9'hb1 == i ? b_177 : _GEN_576;
  assign _GEN_578 = 9'hb2 == i ? b_178 : _GEN_577;
  assign _GEN_579 = 9'hb3 == i ? b_179 : _GEN_578;
  assign _GEN_580 = 9'hb4 == i ? b_180 : _GEN_579;
  assign _GEN_581 = 9'hb5 == i ? b_181 : _GEN_580;
  assign _GEN_582 = 9'hb6 == i ? b_182 : _GEN_581;
  assign _GEN_583 = 9'hb7 == i ? b_183 : _GEN_582;
  assign _GEN_584 = 9'hb8 == i ? b_184 : _GEN_583;
  assign _GEN_585 = 9'hb9 == i ? b_185 : _GEN_584;
  assign _GEN_586 = 9'hba == i ? b_186 : _GEN_585;
  assign _GEN_587 = 9'hbb == i ? b_187 : _GEN_586;
  assign _GEN_588 = 9'hbc == i ? b_188 : _GEN_587;
  assign _GEN_589 = 9'hbd == i ? b_189 : _GEN_588;
  assign _GEN_590 = 9'hbe == i ? b_190 : _GEN_589;
  assign _GEN_591 = 9'hbf == i ? b_191 : _GEN_590;
  assign _GEN_592 = 9'hc0 == i ? b_192 : _GEN_591;
  assign _GEN_593 = 9'hc1 == i ? b_193 : _GEN_592;
  assign _GEN_594 = 9'hc2 == i ? b_194 : _GEN_593;
  assign _GEN_595 = 9'hc3 == i ? b_195 : _GEN_594;
  assign _GEN_596 = 9'hc4 == i ? b_196 : _GEN_595;
  assign _GEN_597 = 9'hc5 == i ? b_197 : _GEN_596;
  assign _GEN_598 = 9'hc6 == i ? b_198 : _GEN_597;
  assign _GEN_599 = 9'hc7 == i ? b_199 : _GEN_598;
  assign _GEN_600 = 9'hc8 == i ? b_200 : _GEN_599;
  assign _GEN_601 = 9'hc9 == i ? b_201 : _GEN_600;
  assign _GEN_602 = 9'hca == i ? b_202 : _GEN_601;
  assign _GEN_603 = 9'hcb == i ? b_203 : _GEN_602;
  assign _GEN_604 = 9'hcc == i ? b_204 : _GEN_603;
  assign _GEN_605 = 9'hcd == i ? b_205 : _GEN_604;
  assign _GEN_606 = 9'hce == i ? b_206 : _GEN_605;
  assign _GEN_607 = 9'hcf == i ? b_207 : _GEN_606;
  assign _GEN_608 = 9'hd0 == i ? b_208 : _GEN_607;
  assign _GEN_609 = 9'hd1 == i ? b_209 : _GEN_608;
  assign _GEN_610 = 9'hd2 == i ? b_210 : _GEN_609;
  assign _GEN_611 = 9'hd3 == i ? b_211 : _GEN_610;
  assign _GEN_612 = 9'hd4 == i ? b_212 : _GEN_611;
  assign _GEN_613 = 9'hd5 == i ? b_213 : _GEN_612;
  assign _GEN_614 = 9'hd6 == i ? b_214 : _GEN_613;
  assign _GEN_615 = 9'hd7 == i ? b_215 : _GEN_614;
  assign _GEN_616 = 9'hd8 == i ? b_216 : _GEN_615;
  assign _GEN_617 = 9'hd9 == i ? b_217 : _GEN_616;
  assign _GEN_618 = 9'hda == i ? b_218 : _GEN_617;
  assign _GEN_619 = 9'hdb == i ? b_219 : _GEN_618;
  assign _GEN_620 = 9'hdc == i ? b_220 : _GEN_619;
  assign _GEN_621 = 9'hdd == i ? b_221 : _GEN_620;
  assign _GEN_622 = 9'hde == i ? b_222 : _GEN_621;
  assign _GEN_623 = 9'hdf == i ? b_223 : _GEN_622;
  assign _GEN_624 = 9'he0 == i ? b_224 : _GEN_623;
  assign _GEN_625 = 9'he1 == i ? b_225 : _GEN_624;
  assign _GEN_626 = 9'he2 == i ? b_226 : _GEN_625;
  assign _GEN_627 = 9'he3 == i ? b_227 : _GEN_626;
  assign _GEN_628 = 9'he4 == i ? b_228 : _GEN_627;
  assign _GEN_629 = 9'he5 == i ? b_229 : _GEN_628;
  assign _GEN_630 = 9'he6 == i ? b_230 : _GEN_629;
  assign _GEN_631 = 9'he7 == i ? b_231 : _GEN_630;
  assign _GEN_632 = 9'he8 == i ? b_232 : _GEN_631;
  assign _GEN_633 = 9'he9 == i ? b_233 : _GEN_632;
  assign _GEN_634 = 9'hea == i ? b_234 : _GEN_633;
  assign _GEN_635 = 9'heb == i ? b_235 : _GEN_634;
  assign _GEN_636 = 9'hec == i ? b_236 : _GEN_635;
  assign _GEN_637 = 9'hed == i ? b_237 : _GEN_636;
  assign _GEN_638 = 9'hee == i ? b_238 : _GEN_637;
  assign _GEN_639 = 9'hef == i ? b_239 : _GEN_638;
  assign _GEN_640 = 9'hf0 == i ? b_240 : _GEN_639;
  assign _GEN_641 = 9'hf1 == i ? b_241 : _GEN_640;
  assign _GEN_642 = 9'hf2 == i ? b_242 : _GEN_641;
  assign _GEN_643 = 9'hf3 == i ? b_243 : _GEN_642;
  assign _GEN_644 = 9'hf4 == i ? b_244 : _GEN_643;
  assign _GEN_645 = 9'hf5 == i ? b_245 : _GEN_644;
  assign _GEN_646 = 9'hf6 == i ? b_246 : _GEN_645;
  assign _GEN_647 = 9'hf7 == i ? b_247 : _GEN_646;
  assign _GEN_648 = 9'hf8 == i ? b_248 : _GEN_647;
  assign _GEN_649 = 9'hf9 == i ? b_249 : _GEN_648;
  assign _GEN_650 = 9'hfa == i ? b_250 : _GEN_649;
  assign _GEN_651 = 9'hfb == i ? b_251 : _GEN_650;
  assign _GEN_652 = 9'hfc == i ? b_252 : _GEN_651;
  assign _GEN_653 = 9'hfd == i ? b_253 : _GEN_652;
  assign _GEN_654 = 9'hfe == i ? b_254 : _GEN_653;
  assign _GEN_655 = 9'hff == i ? b_255 : _GEN_654;
  assign _GEN_656 = 9'h100 == i ? b_256 : _GEN_655;
  assign _GEN_657 = 9'h101 == i ? b_257 : _GEN_656;
  assign _GEN_658 = 9'h102 == i ? b_258 : _GEN_657;
  assign _GEN_659 = 9'h103 == i ? b_259 : _GEN_658;
  assign _GEN_660 = 9'h104 == i ? b_260 : _GEN_659;
  assign _GEN_661 = 9'h105 == i ? b_261 : _GEN_660;
  assign _GEN_662 = 9'h106 == i ? b_262 : _GEN_661;
  assign _GEN_663 = 9'h107 == i ? b_263 : _GEN_662;
  assign _GEN_664 = 9'h108 == i ? b_264 : _GEN_663;
  assign _GEN_665 = 9'h109 == i ? b_265 : _GEN_664;
  assign _GEN_666 = 9'h10a == i ? b_266 : _GEN_665;
  assign _GEN_667 = 9'h10b == i ? b_267 : _GEN_666;
  assign _GEN_668 = 9'h10c == i ? b_268 : _GEN_667;
  assign _GEN_669 = 9'h10d == i ? b_269 : _GEN_668;
  assign _GEN_670 = 9'h10e == i ? b_270 : _GEN_669;
  assign _GEN_671 = 9'h10f == i ? b_271 : _GEN_670;
  assign _GEN_672 = 9'h110 == i ? b_272 : _GEN_671;
  assign _GEN_673 = 9'h111 == i ? b_273 : _GEN_672;
  assign _GEN_674 = 9'h112 == i ? b_274 : _GEN_673;
  assign _GEN_675 = 9'h113 == i ? b_275 : _GEN_674;
  assign _GEN_676 = 9'h114 == i ? b_276 : _GEN_675;
  assign _GEN_677 = 9'h115 == i ? b_277 : _GEN_676;
  assign _GEN_678 = 9'h116 == i ? b_278 : _GEN_677;
  assign _GEN_679 = 9'h117 == i ? b_279 : _GEN_678;
  assign _GEN_680 = 9'h118 == i ? b_280 : _GEN_679;
  assign _GEN_681 = 9'h119 == i ? b_281 : _GEN_680;
  assign _GEN_682 = 9'h11a == i ? b_282 : _GEN_681;
  assign _GEN_683 = 9'h11b == i ? b_283 : _GEN_682;
  assign _GEN_684 = 9'h11c == i ? b_284 : _GEN_683;
  assign _GEN_685 = 9'h11d == i ? b_285 : _GEN_684;
  assign _GEN_686 = 9'h11e == i ? b_286 : _GEN_685;
  assign _GEN_687 = 9'h11f == i ? b_287 : _GEN_686;
  assign _GEN_688 = 9'h120 == i ? b_288 : _GEN_687;
  assign _GEN_689 = 9'h121 == i ? b_289 : _GEN_688;
  assign _GEN_690 = 9'h122 == i ? b_290 : _GEN_689;
  assign _GEN_691 = 9'h123 == i ? b_291 : _GEN_690;
  assign _GEN_692 = 9'h124 == i ? b_292 : _GEN_691;
  assign _GEN_693 = 9'h125 == i ? b_293 : _GEN_692;
  assign _GEN_694 = 9'h126 == i ? b_294 : _GEN_693;
  assign _GEN_695 = 9'h127 == i ? b_295 : _GEN_694;
  assign _GEN_696 = 9'h128 == i ? b_296 : _GEN_695;
  assign _GEN_697 = 9'h129 == i ? b_297 : _GEN_696;
  assign _GEN_698 = 9'h12a == i ? b_298 : _GEN_697;
  assign _GEN_699 = 9'h12b == i ? b_299 : _GEN_698;
  assign _GEN_700 = 9'h12c == i ? b_300 : _GEN_699;
  assign _GEN_701 = 9'h12d == i ? b_301 : _GEN_700;
  assign _GEN_702 = 9'h12e == i ? b_302 : _GEN_701;
  assign _GEN_703 = 9'h12f == i ? b_303 : _GEN_702;
  assign _GEN_704 = 9'h130 == i ? b_304 : _GEN_703;
  assign _GEN_705 = 9'h131 == i ? b_305 : _GEN_704;
  assign _GEN_706 = 9'h132 == i ? b_306 : _GEN_705;
  assign _GEN_707 = 9'h133 == i ? b_307 : _GEN_706;
  assign _GEN_708 = 9'h134 == i ? b_308 : _GEN_707;
  assign _GEN_709 = 9'h135 == i ? b_309 : _GEN_708;
  assign _GEN_710 = 9'h136 == i ? b_310 : _GEN_709;
  assign _GEN_711 = 9'h137 == i ? b_311 : _GEN_710;
  assign _GEN_712 = 9'h138 == i ? b_312 : _GEN_711;
  assign _GEN_713 = 9'h139 == i ? b_313 : _GEN_712;
  assign _GEN_714 = 9'h13a == i ? b_314 : _GEN_713;
  assign _GEN_715 = 9'h13b == i ? b_315 : _GEN_714;
  assign _GEN_716 = 9'h13c == i ? b_316 : _GEN_715;
  assign _GEN_717 = 9'h13d == i ? b_317 : _GEN_716;
  assign _GEN_718 = 9'h13e == i ? b_318 : _GEN_717;
  assign _GEN_719 = 9'h13f == i ? b_319 : _GEN_718;
  assign _GEN_720 = 9'h140 == i ? b_320 : _GEN_719;
  assign _GEN_721 = 9'h141 == i ? b_321 : _GEN_720;
  assign _GEN_722 = 9'h142 == i ? b_322 : _GEN_721;
  assign _GEN_723 = 9'h143 == i ? b_323 : _GEN_722;
  assign _GEN_724 = 9'h144 == i ? b_324 : _GEN_723;
  assign _GEN_725 = 9'h145 == i ? b_325 : _GEN_724;
  assign _GEN_726 = 9'h146 == i ? b_326 : _GEN_725;
  assign _GEN_727 = 9'h147 == i ? b_327 : _GEN_726;
  assign _GEN_728 = 9'h148 == i ? b_328 : _GEN_727;
  assign _GEN_729 = 9'h149 == i ? b_329 : _GEN_728;
  assign _GEN_730 = 9'h14a == i ? b_330 : _GEN_729;
  assign _GEN_731 = 9'h14b == i ? b_331 : _GEN_730;
  assign _GEN_732 = 9'h14c == i ? b_332 : _GEN_731;
  assign _GEN_733 = 9'h14d == i ? b_333 : _GEN_732;
  assign _GEN_734 = 9'h14e == i ? b_334 : _GEN_733;
  assign _GEN_735 = 9'h14f == i ? b_335 : _GEN_734;
  assign _GEN_736 = 9'h150 == i ? b_336 : _GEN_735;
  assign _GEN_737 = 9'h151 == i ? b_337 : _GEN_736;
  assign _GEN_738 = 9'h152 == i ? b_338 : _GEN_737;
  assign _GEN_739 = 9'h153 == i ? b_339 : _GEN_738;
  assign _GEN_740 = 9'h154 == i ? b_340 : _GEN_739;
  assign _GEN_741 = 9'h155 == i ? b_341 : _GEN_740;
  assign _GEN_742 = 9'h156 == i ? b_342 : _GEN_741;
  assign _GEN_743 = 9'h157 == i ? b_343 : _GEN_742;
  assign _GEN_744 = 9'h158 == i ? b_344 : _GEN_743;
  assign _GEN_745 = 9'h159 == i ? b_345 : _GEN_744;
  assign _GEN_746 = 9'h15a == i ? b_346 : _GEN_745;
  assign _GEN_747 = 9'h15b == i ? b_347 : _GEN_746;
  assign _GEN_748 = 9'h15c == i ? b_348 : _GEN_747;
  assign _GEN_749 = 9'h15d == i ? b_349 : _GEN_748;
  assign _GEN_750 = 9'h15e == i ? b_350 : _GEN_749;
  assign _GEN_751 = 9'h15f == i ? b_351 : _GEN_750;
  assign _GEN_752 = 9'h160 == i ? b_352 : _GEN_751;
  assign _GEN_753 = 9'h161 == i ? b_353 : _GEN_752;
  assign _GEN_754 = 9'h162 == i ? b_354 : _GEN_753;
  assign _GEN_755 = 9'h163 == i ? b_355 : _GEN_754;
  assign _GEN_756 = 9'h164 == i ? b_356 : _GEN_755;
  assign _GEN_757 = 9'h165 == i ? b_357 : _GEN_756;
  assign _GEN_758 = 9'h166 == i ? b_358 : _GEN_757;
  assign _GEN_759 = 9'h167 == i ? b_359 : _GEN_758;
  assign _GEN_760 = 9'h168 == i ? b_360 : _GEN_759;
  assign _GEN_761 = 9'h169 == i ? b_361 : _GEN_760;
  assign _GEN_762 = 9'h16a == i ? b_362 : _GEN_761;
  assign _GEN_763 = 9'h16b == i ? b_363 : _GEN_762;
  assign _GEN_764 = 9'h16c == i ? b_364 : _GEN_763;
  assign _GEN_765 = 9'h16d == i ? b_365 : _GEN_764;
  assign _GEN_766 = 9'h16e == i ? b_366 : _GEN_765;
  assign _GEN_767 = 9'h16f == i ? b_367 : _GEN_766;
  assign _GEN_768 = 9'h170 == i ? b_368 : _GEN_767;
  assign _GEN_769 = 9'h171 == i ? b_369 : _GEN_768;
  assign _GEN_770 = 9'h172 == i ? b_370 : _GEN_769;
  assign _GEN_771 = 9'h173 == i ? b_371 : _GEN_770;
  assign _GEN_772 = 9'h174 == i ? b_372 : _GEN_771;
  assign _GEN_773 = 9'h175 == i ? b_373 : _GEN_772;
  assign _GEN_774 = 9'h176 == i ? b_374 : _GEN_773;
  assign _GEN_775 = 9'h177 == i ? b_375 : _GEN_774;
  assign _GEN_776 = 9'h178 == i ? b_376 : _GEN_775;
  assign _GEN_777 = 9'h179 == i ? b_377 : _GEN_776;
  assign _GEN_778 = 9'h17a == i ? b_378 : _GEN_777;
  assign _GEN_779 = 9'h17b == i ? b_379 : _GEN_778;
  assign _GEN_780 = 9'h17c == i ? b_380 : _GEN_779;
  assign _GEN_781 = 9'h17d == i ? b_381 : _GEN_780;
  assign _GEN_782 = 9'h17e == i ? b_382 : _GEN_781;
  assign _GEN_783 = 9'h17f == i ? b_383 : _GEN_782;
  assign _GEN_784 = 9'h180 == i ? b_384 : _GEN_783;
  assign _GEN_785 = 9'h181 == i ? b_385 : _GEN_784;
  assign _GEN_786 = 9'h182 == i ? b_386 : _GEN_785;
  assign _GEN_787 = 9'h183 == i ? b_387 : _GEN_786;
  assign _GEN_788 = 9'h184 == i ? b_388 : _GEN_787;
  assign _GEN_789 = 9'h185 == i ? b_389 : _GEN_788;
  assign _GEN_790 = 9'h186 == i ? b_390 : _GEN_789;
  assign _GEN_791 = 9'h187 == i ? b_391 : _GEN_790;
  assign _GEN_792 = 9'h188 == i ? b_392 : _GEN_791;
  assign _GEN_793 = 9'h189 == i ? b_393 : _GEN_792;
  assign _GEN_794 = 9'h18a == i ? b_394 : _GEN_793;
  assign _GEN_795 = 9'h18b == i ? b_395 : _GEN_794;
  assign _GEN_796 = 9'h18c == i ? b_396 : _GEN_795;
  assign _GEN_797 = 9'h18d == i ? b_397 : _GEN_796;
  assign _GEN_798 = 9'h18e == i ? b_398 : _GEN_797;
  assign _GEN_799 = 9'h18f == i ? b_399 : _GEN_798;
  assign _T_800 = _GEN_399 * _GEN_799;
  assign _T_801 = sum + _T_800;
  assign _T_802 = i + 9'h1;
  assign _GEN_800 = _T_804 ? _T_802 : 10'h0;
  assign _GEN_801 = _T_804 ? _T_801 : 33'h0;
  assign _GEN_802 = _T_803 ? 10'h0 : _GEN_800;
  assign _GEN_804 = _T_803 ? sum : 32'h0;
  assign _GEN_805 = _T_803 ? 33'h0 : _GEN_801;
  assign _GEN_806 = io_rdy ? _T_801 : _GEN_805;
  assign _GEN_807 = io_rdy ? _T_802 : _GEN_802;
  assign io_q = io_rdy ? 32'h0 : _GEN_804;
  assign io_v = io_rdy ? 1'h0 : _T_803;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sum = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  i = _RAND_1[8:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      sum <= 32'h0;
    end else begin
      sum <= _GEN_806[31:0];
    end
    if (reset) begin
      i <= 9'h0;
    end else begin
      i <= _GEN_807[8:0];
    end
  end
endmodule
module Node_102(
  input           clock,
  input           reset,
  input  [6399:0] io_d_in,
  input  [6399:0] io_w,
  input           io_rdy,
  input  [15:0]   io_bias,
  output [15:0]   io_d_out,
  output          io_v
);
  wire  muladdc_clock;
  wire  muladdc_reset;
  wire [6399:0] muladdc_io_a;
  wire [6399:0] muladdc_io_b;
  wire  muladdc_io_rdy;
  wire [31:0] muladdc_io_q;
  wire  muladdc_io_v;
  wire [31:0] act_io_q;
  wire [15:0] act_io_bias;
  wire  act_io_v_in;
  wire [15:0] act_io_d;
  wire  act_io_v_out;
  Mac_102 muladdc (
    .clock(muladdc_clock),
    .reset(muladdc_reset),
    .io_a(muladdc_io_a),
    .io_b(muladdc_io_b),
    .io_rdy(muladdc_io_rdy),
    .io_q(muladdc_io_q),
    .io_v(muladdc_io_v)
  );
  ReLU act (
    .io_q(act_io_q),
    .io_bias(act_io_bias),
    .io_v_in(act_io_v_in),
    .io_d(act_io_d),
    .io_v_out(act_io_v_out)
  );
  assign io_d_out = act_io_d;
  assign io_v = act_io_v_out;
  assign muladdc_clock = clock;
  assign muladdc_reset = reset;
  assign muladdc_io_a = io_d_in;
  assign muladdc_io_b = io_w;
  assign muladdc_io_rdy = io_rdy;
  assign act_io_q = muladdc_io_q;
  assign act_io_bias = io_bias;
  assign act_io_v_in = muladdc_io_v;
endmodule
module FC1(
  input           clock,
  input           reset,
  input  [15:0]   io_d_in_0,
  input  [15:0]   io_d_in_1,
  input  [15:0]   io_d_in_2,
  input  [15:0]   io_d_in_3,
  input  [15:0]   io_d_in_4,
  input  [15:0]   io_d_in_5,
  input  [15:0]   io_d_in_6,
  input  [15:0]   io_d_in_7,
  input  [15:0]   io_d_in_8,
  input  [15:0]   io_d_in_9,
  input  [15:0]   io_d_in_10,
  input  [15:0]   io_d_in_11,
  input  [15:0]   io_d_in_12,
  input  [15:0]   io_d_in_13,
  input  [15:0]   io_d_in_14,
  input  [15:0]   io_d_in_15,
  input  [3199:0] io_wa_in,
  input  [3199:0] io_wb_in,
  input  [15:0]   io_bias,
  input           io_rdy,
  input           io_done,
  output [15:0]   io_d_out,
  output          io_v
);
  wire  _T_1_clock;
  wire  _T_1_reset;
  wire [15:0] _T_1_io_d_in;
  wire  _T_1_io_en;
  wire [399:0] _T_1_io_d_out;
  wire  _T_2_clock;
  wire  _T_2_reset;
  wire [15:0] _T_2_io_d_in;
  wire  _T_2_io_en;
  wire [399:0] _T_2_io_d_out;
  wire  _T_4_clock;
  wire  _T_4_reset;
  wire [15:0] _T_4_io_d_in;
  wire  _T_4_io_en;
  wire [399:0] _T_4_io_d_out;
  wire  _T_5_clock;
  wire  _T_5_reset;
  wire [15:0] _T_5_io_d_in;
  wire  _T_5_io_en;
  wire [399:0] _T_5_io_d_out;
  wire  _T_8_clock;
  wire  _T_8_reset;
  wire [15:0] _T_8_io_d_in;
  wire  _T_8_io_en;
  wire [399:0] _T_8_io_d_out;
  wire  _T_9_clock;
  wire  _T_9_reset;
  wire [15:0] _T_9_io_d_in;
  wire  _T_9_io_en;
  wire [399:0] _T_9_io_d_out;
  wire  _T_11_clock;
  wire  _T_11_reset;
  wire [15:0] _T_11_io_d_in;
  wire  _T_11_io_en;
  wire [399:0] _T_11_io_d_out;
  wire  _T_12_clock;
  wire  _T_12_reset;
  wire [15:0] _T_12_io_d_in;
  wire  _T_12_io_en;
  wire [399:0] _T_12_io_d_out;
  wire  _T_16_clock;
  wire  _T_16_reset;
  wire [15:0] _T_16_io_d_in;
  wire  _T_16_io_en;
  wire [399:0] _T_16_io_d_out;
  wire  _T_17_clock;
  wire  _T_17_reset;
  wire [15:0] _T_17_io_d_in;
  wire  _T_17_io_en;
  wire [399:0] _T_17_io_d_out;
  wire  _T_19_clock;
  wire  _T_19_reset;
  wire [15:0] _T_19_io_d_in;
  wire  _T_19_io_en;
  wire [399:0] _T_19_io_d_out;
  wire  _T_20_clock;
  wire  _T_20_reset;
  wire [15:0] _T_20_io_d_in;
  wire  _T_20_io_en;
  wire [399:0] _T_20_io_d_out;
  wire  _T_23_clock;
  wire  _T_23_reset;
  wire [15:0] _T_23_io_d_in;
  wire  _T_23_io_en;
  wire [399:0] _T_23_io_d_out;
  wire  _T_24_clock;
  wire  _T_24_reset;
  wire [15:0] _T_24_io_d_in;
  wire  _T_24_io_en;
  wire [399:0] _T_24_io_d_out;
  wire  _T_26_clock;
  wire  _T_26_reset;
  wire [15:0] _T_26_io_d_in;
  wire  _T_26_io_en;
  wire [399:0] _T_26_io_d_out;
  wire  _T_27_clock;
  wire  _T_27_reset;
  wire [15:0] _T_27_io_d_in;
  wire  _T_27_io_en;
  wire [399:0] _T_27_io_d_out;
  wire  conv_node_clock;
  wire  conv_node_reset;
  wire [6399:0] conv_node_io_d_in;
  wire [6399:0] conv_node_io_w;
  wire  conv_node_io_rdy;
  wire [15:0] conv_node_io_bias;
  wire [15:0] conv_node_io_d_out;
  wire  conv_node_io_v;
  reg [6399:0] din;
  reg [6399:0] _RAND_0;
  reg  first_rdy;
  reg [31:0] _RAND_1;
  reg [15:0] channel_counter;
  reg [31:0] _RAND_2;
  wire  _T;
  wire [3199:0] _T_30;
  wire [6399:0] _T_31;
  wire [16:0] _T_32;
  wire [16:0] _GEN_0;
  wire [16:0] _GEN_1;
  reg  is_done;
  reg [31:0] _RAND_3;
  wire  _GEN_4;
  reg  rdy;
  reg [31:0] _RAND_4;
  wire  _T_34;
  ShiftRegister _T_1 (
    .clock(_T_1_clock),
    .reset(_T_1_reset),
    .io_d_in(_T_1_io_d_in),
    .io_en(_T_1_io_en),
    .io_d_out(_T_1_io_d_out)
  );
  ShiftRegister _T_2 (
    .clock(_T_2_clock),
    .reset(_T_2_reset),
    .io_d_in(_T_2_io_d_in),
    .io_en(_T_2_io_en),
    .io_d_out(_T_2_io_d_out)
  );
  ShiftRegister _T_4 (
    .clock(_T_4_clock),
    .reset(_T_4_reset),
    .io_d_in(_T_4_io_d_in),
    .io_en(_T_4_io_en),
    .io_d_out(_T_4_io_d_out)
  );
  ShiftRegister _T_5 (
    .clock(_T_5_clock),
    .reset(_T_5_reset),
    .io_d_in(_T_5_io_d_in),
    .io_en(_T_5_io_en),
    .io_d_out(_T_5_io_d_out)
  );
  ShiftRegister _T_8 (
    .clock(_T_8_clock),
    .reset(_T_8_reset),
    .io_d_in(_T_8_io_d_in),
    .io_en(_T_8_io_en),
    .io_d_out(_T_8_io_d_out)
  );
  ShiftRegister _T_9 (
    .clock(_T_9_clock),
    .reset(_T_9_reset),
    .io_d_in(_T_9_io_d_in),
    .io_en(_T_9_io_en),
    .io_d_out(_T_9_io_d_out)
  );
  ShiftRegister _T_11 (
    .clock(_T_11_clock),
    .reset(_T_11_reset),
    .io_d_in(_T_11_io_d_in),
    .io_en(_T_11_io_en),
    .io_d_out(_T_11_io_d_out)
  );
  ShiftRegister _T_12 (
    .clock(_T_12_clock),
    .reset(_T_12_reset),
    .io_d_in(_T_12_io_d_in),
    .io_en(_T_12_io_en),
    .io_d_out(_T_12_io_d_out)
  );
  ShiftRegister _T_16 (
    .clock(_T_16_clock),
    .reset(_T_16_reset),
    .io_d_in(_T_16_io_d_in),
    .io_en(_T_16_io_en),
    .io_d_out(_T_16_io_d_out)
  );
  ShiftRegister _T_17 (
    .clock(_T_17_clock),
    .reset(_T_17_reset),
    .io_d_in(_T_17_io_d_in),
    .io_en(_T_17_io_en),
    .io_d_out(_T_17_io_d_out)
  );
  ShiftRegister _T_19 (
    .clock(_T_19_clock),
    .reset(_T_19_reset),
    .io_d_in(_T_19_io_d_in),
    .io_en(_T_19_io_en),
    .io_d_out(_T_19_io_d_out)
  );
  ShiftRegister _T_20 (
    .clock(_T_20_clock),
    .reset(_T_20_reset),
    .io_d_in(_T_20_io_d_in),
    .io_en(_T_20_io_en),
    .io_d_out(_T_20_io_d_out)
  );
  ShiftRegister _T_23 (
    .clock(_T_23_clock),
    .reset(_T_23_reset),
    .io_d_in(_T_23_io_d_in),
    .io_en(_T_23_io_en),
    .io_d_out(_T_23_io_d_out)
  );
  ShiftRegister _T_24 (
    .clock(_T_24_clock),
    .reset(_T_24_reset),
    .io_d_in(_T_24_io_d_in),
    .io_en(_T_24_io_en),
    .io_d_out(_T_24_io_d_out)
  );
  ShiftRegister _T_26 (
    .clock(_T_26_clock),
    .reset(_T_26_reset),
    .io_d_in(_T_26_io_d_in),
    .io_en(_T_26_io_en),
    .io_d_out(_T_26_io_d_out)
  );
  ShiftRegister _T_27 (
    .clock(_T_27_clock),
    .reset(_T_27_reset),
    .io_d_in(_T_27_io_d_in),
    .io_en(_T_27_io_en),
    .io_d_out(_T_27_io_d_out)
  );
  Node_102 conv_node (
    .clock(conv_node_clock),
    .reset(conv_node_reset),
    .io_d_in(conv_node_io_d_in),
    .io_w(conv_node_io_w),
    .io_rdy(conv_node_io_rdy),
    .io_bias(conv_node_io_bias),
    .io_d_out(conv_node_io_d_out),
    .io_v(conv_node_io_v)
  );
  assign _T = channel_counter == 16'h19;
  assign _T_30 = {_T_16_io_d_out,_T_17_io_d_out,_T_19_io_d_out,_T_20_io_d_out,_T_23_io_d_out,_T_24_io_d_out,_T_26_io_d_out,_T_27_io_d_out};
  assign _T_31 = {_T_1_io_d_out,_T_2_io_d_out,_T_4_io_d_out,_T_5_io_d_out,_T_8_io_d_out,_T_9_io_d_out,_T_11_io_d_out,_T_12_io_d_out,_T_30};
  assign _T_32 = channel_counter + 16'h1;
  assign _GEN_0 = io_rdy ? _T_32 : {{1'd0}, channel_counter};
  assign _GEN_1 = _T ? 17'h0 : _GEN_0;
  assign _GEN_4 = io_done | is_done;
  assign _T_34 = first_rdy | conv_node_io_v;
  assign io_d_out = conv_node_io_d_out;
  assign io_v = conv_node_io_v;
  assign _T_1_clock = clock;
  assign _T_1_reset = reset;
  assign _T_1_io_d_in = io_d_in_0;
  assign _T_1_io_en = io_rdy;
  assign _T_2_clock = clock;
  assign _T_2_reset = reset;
  assign _T_2_io_d_in = io_d_in_1;
  assign _T_2_io_en = io_rdy;
  assign _T_4_clock = clock;
  assign _T_4_reset = reset;
  assign _T_4_io_d_in = io_d_in_2;
  assign _T_4_io_en = io_rdy;
  assign _T_5_clock = clock;
  assign _T_5_reset = reset;
  assign _T_5_io_d_in = io_d_in_3;
  assign _T_5_io_en = io_rdy;
  assign _T_8_clock = clock;
  assign _T_8_reset = reset;
  assign _T_8_io_d_in = io_d_in_4;
  assign _T_8_io_en = io_rdy;
  assign _T_9_clock = clock;
  assign _T_9_reset = reset;
  assign _T_9_io_d_in = io_d_in_5;
  assign _T_9_io_en = io_rdy;
  assign _T_11_clock = clock;
  assign _T_11_reset = reset;
  assign _T_11_io_d_in = io_d_in_6;
  assign _T_11_io_en = io_rdy;
  assign _T_12_clock = clock;
  assign _T_12_reset = reset;
  assign _T_12_io_d_in = io_d_in_7;
  assign _T_12_io_en = io_rdy;
  assign _T_16_clock = clock;
  assign _T_16_reset = reset;
  assign _T_16_io_d_in = io_d_in_8;
  assign _T_16_io_en = io_rdy;
  assign _T_17_clock = clock;
  assign _T_17_reset = reset;
  assign _T_17_io_d_in = io_d_in_9;
  assign _T_17_io_en = io_rdy;
  assign _T_19_clock = clock;
  assign _T_19_reset = reset;
  assign _T_19_io_d_in = io_d_in_10;
  assign _T_19_io_en = io_rdy;
  assign _T_20_clock = clock;
  assign _T_20_reset = reset;
  assign _T_20_io_d_in = io_d_in_11;
  assign _T_20_io_en = io_rdy;
  assign _T_23_clock = clock;
  assign _T_23_reset = reset;
  assign _T_23_io_d_in = io_d_in_12;
  assign _T_23_io_en = io_rdy;
  assign _T_24_clock = clock;
  assign _T_24_reset = reset;
  assign _T_24_io_d_in = io_d_in_13;
  assign _T_24_io_en = io_rdy;
  assign _T_26_clock = clock;
  assign _T_26_reset = reset;
  assign _T_26_io_d_in = io_d_in_14;
  assign _T_26_io_en = io_rdy;
  assign _T_27_clock = clock;
  assign _T_27_reset = reset;
  assign _T_27_io_d_in = io_d_in_15;
  assign _T_27_io_en = io_rdy;
  assign conv_node_clock = clock;
  assign conv_node_reset = reset;
  assign conv_node_io_d_in = din;
  assign conv_node_io_w = {io_wa_in,io_wb_in};
  assign conv_node_io_rdy = rdy;
  assign conv_node_io_bias = io_bias;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {200{`RANDOM}};
  din = _RAND_0[6399:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  first_rdy = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  channel_counter = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  is_done = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  rdy = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      din <= 'h0;
    end else if (_T) begin
      din <= _T_31;
    end
    if (reset) begin
      first_rdy <= 1'h0;
    end else begin
      first_rdy <= _T;
    end
    if (reset) begin
      channel_counter <= 16'h0;
    end else begin
      channel_counter <= _GEN_1[15:0];
    end
    if (reset) begin
      is_done <= 1'h0;
    end else begin
      is_done <= _GEN_4;
    end
    if (reset) begin
      rdy <= 1'h0;
    end else if (is_done) begin
      rdy <= 1'h0;
    end else begin
      rdy <= _T_34;
    end
  end
endmodule
module ShiftRegister_22(
  input           clock,
  input           reset,
  input  [15:0]   io_d_in,
  input           io_en,
  output [1919:0] io_d_out
);
  reg [15:0] _T;
  reg [31:0] _RAND_0;
  reg [15:0] _T_1;
  reg [31:0] _RAND_1;
  reg [15:0] _T_2;
  reg [31:0] _RAND_2;
  reg [15:0] _T_3;
  reg [31:0] _RAND_3;
  reg [15:0] _T_4;
  reg [31:0] _RAND_4;
  reg [15:0] _T_5;
  reg [31:0] _RAND_5;
  reg [15:0] _T_6;
  reg [31:0] _RAND_6;
  reg [15:0] _T_7;
  reg [31:0] _RAND_7;
  reg [15:0] _T_8;
  reg [31:0] _RAND_8;
  reg [15:0] _T_9;
  reg [31:0] _RAND_9;
  reg [15:0] _T_10;
  reg [31:0] _RAND_10;
  reg [15:0] _T_11;
  reg [31:0] _RAND_11;
  reg [15:0] _T_12;
  reg [31:0] _RAND_12;
  reg [15:0] _T_13;
  reg [31:0] _RAND_13;
  reg [15:0] _T_14;
  reg [31:0] _RAND_14;
  reg [15:0] _T_15;
  reg [31:0] _RAND_15;
  reg [15:0] _T_16;
  reg [31:0] _RAND_16;
  reg [15:0] _T_17;
  reg [31:0] _RAND_17;
  reg [15:0] _T_18;
  reg [31:0] _RAND_18;
  reg [15:0] _T_19;
  reg [31:0] _RAND_19;
  reg [15:0] _T_20;
  reg [31:0] _RAND_20;
  reg [15:0] _T_21;
  reg [31:0] _RAND_21;
  reg [15:0] _T_22;
  reg [31:0] _RAND_22;
  reg [15:0] _T_23;
  reg [31:0] _RAND_23;
  reg [15:0] _T_24;
  reg [31:0] _RAND_24;
  reg [15:0] _T_25;
  reg [31:0] _RAND_25;
  reg [15:0] _T_26;
  reg [31:0] _RAND_26;
  reg [15:0] _T_27;
  reg [31:0] _RAND_27;
  reg [15:0] _T_28;
  reg [31:0] _RAND_28;
  reg [15:0] _T_29;
  reg [31:0] _RAND_29;
  reg [15:0] _T_30;
  reg [31:0] _RAND_30;
  reg [15:0] _T_31;
  reg [31:0] _RAND_31;
  reg [15:0] _T_32;
  reg [31:0] _RAND_32;
  reg [15:0] _T_33;
  reg [31:0] _RAND_33;
  reg [15:0] _T_34;
  reg [31:0] _RAND_34;
  reg [15:0] _T_35;
  reg [31:0] _RAND_35;
  reg [15:0] _T_36;
  reg [31:0] _RAND_36;
  reg [15:0] _T_37;
  reg [31:0] _RAND_37;
  reg [15:0] _T_38;
  reg [31:0] _RAND_38;
  reg [15:0] _T_39;
  reg [31:0] _RAND_39;
  reg [15:0] _T_40;
  reg [31:0] _RAND_40;
  reg [15:0] _T_41;
  reg [31:0] _RAND_41;
  reg [15:0] _T_42;
  reg [31:0] _RAND_42;
  reg [15:0] _T_43;
  reg [31:0] _RAND_43;
  reg [15:0] _T_44;
  reg [31:0] _RAND_44;
  reg [15:0] _T_45;
  reg [31:0] _RAND_45;
  reg [15:0] _T_46;
  reg [31:0] _RAND_46;
  reg [15:0] _T_47;
  reg [31:0] _RAND_47;
  reg [15:0] _T_48;
  reg [31:0] _RAND_48;
  reg [15:0] _T_49;
  reg [31:0] _RAND_49;
  reg [15:0] _T_50;
  reg [31:0] _RAND_50;
  reg [15:0] _T_51;
  reg [31:0] _RAND_51;
  reg [15:0] _T_52;
  reg [31:0] _RAND_52;
  reg [15:0] _T_53;
  reg [31:0] _RAND_53;
  reg [15:0] _T_54;
  reg [31:0] _RAND_54;
  reg [15:0] _T_55;
  reg [31:0] _RAND_55;
  reg [15:0] _T_56;
  reg [31:0] _RAND_56;
  reg [15:0] _T_57;
  reg [31:0] _RAND_57;
  reg [15:0] _T_58;
  reg [31:0] _RAND_58;
  reg [15:0] _T_59;
  reg [31:0] _RAND_59;
  reg [15:0] _T_60;
  reg [31:0] _RAND_60;
  reg [15:0] _T_61;
  reg [31:0] _RAND_61;
  reg [15:0] _T_62;
  reg [31:0] _RAND_62;
  reg [15:0] _T_63;
  reg [31:0] _RAND_63;
  reg [15:0] _T_64;
  reg [31:0] _RAND_64;
  reg [15:0] _T_65;
  reg [31:0] _RAND_65;
  reg [15:0] _T_66;
  reg [31:0] _RAND_66;
  reg [15:0] _T_67;
  reg [31:0] _RAND_67;
  reg [15:0] _T_68;
  reg [31:0] _RAND_68;
  reg [15:0] _T_69;
  reg [31:0] _RAND_69;
  reg [15:0] _T_70;
  reg [31:0] _RAND_70;
  reg [15:0] _T_71;
  reg [31:0] _RAND_71;
  reg [15:0] _T_72;
  reg [31:0] _RAND_72;
  reg [15:0] _T_73;
  reg [31:0] _RAND_73;
  reg [15:0] _T_74;
  reg [31:0] _RAND_74;
  reg [15:0] _T_75;
  reg [31:0] _RAND_75;
  reg [15:0] _T_76;
  reg [31:0] _RAND_76;
  reg [15:0] _T_77;
  reg [31:0] _RAND_77;
  reg [15:0] _T_78;
  reg [31:0] _RAND_78;
  reg [15:0] _T_79;
  reg [31:0] _RAND_79;
  reg [15:0] _T_80;
  reg [31:0] _RAND_80;
  reg [15:0] _T_81;
  reg [31:0] _RAND_81;
  reg [15:0] _T_82;
  reg [31:0] _RAND_82;
  reg [15:0] _T_83;
  reg [31:0] _RAND_83;
  reg [15:0] _T_84;
  reg [31:0] _RAND_84;
  reg [15:0] _T_85;
  reg [31:0] _RAND_85;
  reg [15:0] _T_86;
  reg [31:0] _RAND_86;
  reg [15:0] _T_87;
  reg [31:0] _RAND_87;
  reg [15:0] _T_88;
  reg [31:0] _RAND_88;
  reg [15:0] _T_89;
  reg [31:0] _RAND_89;
  reg [15:0] _T_90;
  reg [31:0] _RAND_90;
  reg [15:0] _T_91;
  reg [31:0] _RAND_91;
  reg [15:0] _T_92;
  reg [31:0] _RAND_92;
  reg [15:0] _T_93;
  reg [31:0] _RAND_93;
  reg [15:0] _T_94;
  reg [31:0] _RAND_94;
  reg [15:0] _T_95;
  reg [31:0] _RAND_95;
  reg [15:0] _T_96;
  reg [31:0] _RAND_96;
  reg [15:0] _T_97;
  reg [31:0] _RAND_97;
  reg [15:0] _T_98;
  reg [31:0] _RAND_98;
  reg [15:0] _T_99;
  reg [31:0] _RAND_99;
  reg [15:0] _T_100;
  reg [31:0] _RAND_100;
  reg [15:0] _T_101;
  reg [31:0] _RAND_101;
  reg [15:0] _T_102;
  reg [31:0] _RAND_102;
  reg [15:0] _T_103;
  reg [31:0] _RAND_103;
  reg [15:0] _T_104;
  reg [31:0] _RAND_104;
  reg [15:0] _T_105;
  reg [31:0] _RAND_105;
  reg [15:0] _T_106;
  reg [31:0] _RAND_106;
  reg [15:0] _T_107;
  reg [31:0] _RAND_107;
  reg [15:0] _T_108;
  reg [31:0] _RAND_108;
  reg [15:0] _T_109;
  reg [31:0] _RAND_109;
  reg [15:0] _T_110;
  reg [31:0] _RAND_110;
  reg [15:0] _T_111;
  reg [31:0] _RAND_111;
  reg [15:0] _T_112;
  reg [31:0] _RAND_112;
  reg [15:0] _T_113;
  reg [31:0] _RAND_113;
  reg [15:0] _T_114;
  reg [31:0] _RAND_114;
  reg [15:0] _T_115;
  reg [31:0] _RAND_115;
  reg [15:0] _T_116;
  reg [31:0] _RAND_116;
  reg [15:0] _T_117;
  reg [31:0] _RAND_117;
  reg [15:0] _T_118;
  reg [31:0] _RAND_118;
  reg [15:0] _T_119;
  reg [31:0] _RAND_119;
  wire [127:0] _T_132;
  wire [127:0] _T_146;
  wire [239:0] _T_147;
  wire [127:0] _T_161;
  wire [127:0] _T_175;
  wire [239:0] _T_176;
  wire [479:0] _T_177;
  wire [959:0] _T_178;
  wire [127:0] _T_191;
  wire [127:0] _T_205;
  wire [239:0] _T_206;
  wire [127:0] _T_220;
  wire [127:0] _T_234;
  wire [239:0] _T_235;
  wire [479:0] _T_236;
  wire [959:0] _T_237;
  assign _T_132 = {_T_7,_T_8,_T_9,_T_10,_T_11,_T_12,_T_13,_T_14};
  assign _T_146 = {_T_22,_T_23,_T_24,_T_25,_T_26,_T_27,_T_28,_T_29};
  assign _T_147 = {_T_15,_T_16,_T_17,_T_18,_T_19,_T_20,_T_21,_T_146};
  assign _T_161 = {_T_37,_T_38,_T_39,_T_40,_T_41,_T_42,_T_43,_T_44};
  assign _T_175 = {_T_52,_T_53,_T_54,_T_55,_T_56,_T_57,_T_58,_T_59};
  assign _T_176 = {_T_45,_T_46,_T_47,_T_48,_T_49,_T_50,_T_51,_T_175};
  assign _T_177 = {_T_30,_T_31,_T_32,_T_33,_T_34,_T_35,_T_36,_T_161,_T_176};
  assign _T_178 = {_T,_T_1,_T_2,_T_3,_T_4,_T_5,_T_6,_T_132,_T_147,_T_177};
  assign _T_191 = {_T_67,_T_68,_T_69,_T_70,_T_71,_T_72,_T_73,_T_74};
  assign _T_205 = {_T_82,_T_83,_T_84,_T_85,_T_86,_T_87,_T_88,_T_89};
  assign _T_206 = {_T_75,_T_76,_T_77,_T_78,_T_79,_T_80,_T_81,_T_205};
  assign _T_220 = {_T_97,_T_98,_T_99,_T_100,_T_101,_T_102,_T_103,_T_104};
  assign _T_234 = {_T_112,_T_113,_T_114,_T_115,_T_116,_T_117,_T_118,_T_119};
  assign _T_235 = {_T_105,_T_106,_T_107,_T_108,_T_109,_T_110,_T_111,_T_234};
  assign _T_236 = {_T_90,_T_91,_T_92,_T_93,_T_94,_T_95,_T_96,_T_220,_T_235};
  assign _T_237 = {_T_60,_T_61,_T_62,_T_63,_T_64,_T_65,_T_66,_T_191,_T_206,_T_236};
  assign io_d_out = {_T_178,_T_237};
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_6 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_7 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_8 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_9 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_10 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_11 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_12 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_13 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_14 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_15 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_16 = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_17 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_18 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_19 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_20 = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_21 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_22 = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_23 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_24 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_25 = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_26 = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_27 = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_28 = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_29 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_30 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_31 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_32 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_33 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_34 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_35 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_36 = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_37 = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_38 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_39 = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_40 = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_41 = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_42 = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_43 = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_44 = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_45 = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_46 = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_47 = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_48 = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_49 = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_50 = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_51 = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_52 = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_53 = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_54 = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_55 = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_56 = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_57 = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_58 = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_59 = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_60 = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_61 = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_62 = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_63 = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_64 = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_65 = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_66 = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_67 = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_68 = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_69 = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_70 = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_71 = _RAND_71[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_72 = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_73 = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_74 = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_75 = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_76 = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_77 = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_78 = _RAND_78[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_79 = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_80 = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_81 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_82 = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_83 = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_84 = _RAND_84[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_85 = _RAND_85[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_86 = _RAND_86[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_87 = _RAND_87[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_88 = _RAND_88[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_89 = _RAND_89[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_90 = _RAND_90[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_91 = _RAND_91[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_92 = _RAND_92[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_93 = _RAND_93[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_94 = _RAND_94[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_95 = _RAND_95[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_96 = _RAND_96[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_97 = _RAND_97[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_98 = _RAND_98[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_99 = _RAND_99[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_100 = _RAND_100[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_101 = _RAND_101[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_102 = _RAND_102[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_103 = _RAND_103[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_104 = _RAND_104[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_105 = _RAND_105[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_106 = _RAND_106[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_107 = _RAND_107[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_108 = _RAND_108[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_109 = _RAND_109[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_110 = _RAND_110[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_111 = _RAND_111[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_112 = _RAND_112[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_113 = _RAND_113[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_114 = _RAND_114[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_115 = _RAND_115[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_116 = _RAND_116[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_117 = _RAND_117[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_118 = _RAND_118[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_119 = _RAND_119[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T <= 16'h0;
    end else if (io_en) begin
      _T <= io_d_in;
    end
    if (reset) begin
      _T_1 <= 16'h0;
    end else if (io_en) begin
      _T_1 <= _T;
    end
    if (reset) begin
      _T_2 <= 16'h0;
    end else if (io_en) begin
      _T_2 <= _T_1;
    end
    if (reset) begin
      _T_3 <= 16'h0;
    end else if (io_en) begin
      _T_3 <= _T_2;
    end
    if (reset) begin
      _T_4 <= 16'h0;
    end else if (io_en) begin
      _T_4 <= _T_3;
    end
    if (reset) begin
      _T_5 <= 16'h0;
    end else if (io_en) begin
      _T_5 <= _T_4;
    end
    if (reset) begin
      _T_6 <= 16'h0;
    end else if (io_en) begin
      _T_6 <= _T_5;
    end
    if (reset) begin
      _T_7 <= 16'h0;
    end else if (io_en) begin
      _T_7 <= _T_6;
    end
    if (reset) begin
      _T_8 <= 16'h0;
    end else if (io_en) begin
      _T_8 <= _T_7;
    end
    if (reset) begin
      _T_9 <= 16'h0;
    end else if (io_en) begin
      _T_9 <= _T_8;
    end
    if (reset) begin
      _T_10 <= 16'h0;
    end else if (io_en) begin
      _T_10 <= _T_9;
    end
    if (reset) begin
      _T_11 <= 16'h0;
    end else if (io_en) begin
      _T_11 <= _T_10;
    end
    if (reset) begin
      _T_12 <= 16'h0;
    end else if (io_en) begin
      _T_12 <= _T_11;
    end
    if (reset) begin
      _T_13 <= 16'h0;
    end else if (io_en) begin
      _T_13 <= _T_12;
    end
    if (reset) begin
      _T_14 <= 16'h0;
    end else if (io_en) begin
      _T_14 <= _T_13;
    end
    if (reset) begin
      _T_15 <= 16'h0;
    end else if (io_en) begin
      _T_15 <= _T_14;
    end
    if (reset) begin
      _T_16 <= 16'h0;
    end else if (io_en) begin
      _T_16 <= _T_15;
    end
    if (reset) begin
      _T_17 <= 16'h0;
    end else if (io_en) begin
      _T_17 <= _T_16;
    end
    if (reset) begin
      _T_18 <= 16'h0;
    end else if (io_en) begin
      _T_18 <= _T_17;
    end
    if (reset) begin
      _T_19 <= 16'h0;
    end else if (io_en) begin
      _T_19 <= _T_18;
    end
    if (reset) begin
      _T_20 <= 16'h0;
    end else if (io_en) begin
      _T_20 <= _T_19;
    end
    if (reset) begin
      _T_21 <= 16'h0;
    end else if (io_en) begin
      _T_21 <= _T_20;
    end
    if (reset) begin
      _T_22 <= 16'h0;
    end else if (io_en) begin
      _T_22 <= _T_21;
    end
    if (reset) begin
      _T_23 <= 16'h0;
    end else if (io_en) begin
      _T_23 <= _T_22;
    end
    if (reset) begin
      _T_24 <= 16'h0;
    end else if (io_en) begin
      _T_24 <= _T_23;
    end
    if (reset) begin
      _T_25 <= 16'h0;
    end else if (io_en) begin
      _T_25 <= _T_24;
    end
    if (reset) begin
      _T_26 <= 16'h0;
    end else if (io_en) begin
      _T_26 <= _T_25;
    end
    if (reset) begin
      _T_27 <= 16'h0;
    end else if (io_en) begin
      _T_27 <= _T_26;
    end
    if (reset) begin
      _T_28 <= 16'h0;
    end else if (io_en) begin
      _T_28 <= _T_27;
    end
    if (reset) begin
      _T_29 <= 16'h0;
    end else if (io_en) begin
      _T_29 <= _T_28;
    end
    if (reset) begin
      _T_30 <= 16'h0;
    end else if (io_en) begin
      _T_30 <= _T_29;
    end
    if (reset) begin
      _T_31 <= 16'h0;
    end else if (io_en) begin
      _T_31 <= _T_30;
    end
    if (reset) begin
      _T_32 <= 16'h0;
    end else if (io_en) begin
      _T_32 <= _T_31;
    end
    if (reset) begin
      _T_33 <= 16'h0;
    end else if (io_en) begin
      _T_33 <= _T_32;
    end
    if (reset) begin
      _T_34 <= 16'h0;
    end else if (io_en) begin
      _T_34 <= _T_33;
    end
    if (reset) begin
      _T_35 <= 16'h0;
    end else if (io_en) begin
      _T_35 <= _T_34;
    end
    if (reset) begin
      _T_36 <= 16'h0;
    end else if (io_en) begin
      _T_36 <= _T_35;
    end
    if (reset) begin
      _T_37 <= 16'h0;
    end else if (io_en) begin
      _T_37 <= _T_36;
    end
    if (reset) begin
      _T_38 <= 16'h0;
    end else if (io_en) begin
      _T_38 <= _T_37;
    end
    if (reset) begin
      _T_39 <= 16'h0;
    end else if (io_en) begin
      _T_39 <= _T_38;
    end
    if (reset) begin
      _T_40 <= 16'h0;
    end else if (io_en) begin
      _T_40 <= _T_39;
    end
    if (reset) begin
      _T_41 <= 16'h0;
    end else if (io_en) begin
      _T_41 <= _T_40;
    end
    if (reset) begin
      _T_42 <= 16'h0;
    end else if (io_en) begin
      _T_42 <= _T_41;
    end
    if (reset) begin
      _T_43 <= 16'h0;
    end else if (io_en) begin
      _T_43 <= _T_42;
    end
    if (reset) begin
      _T_44 <= 16'h0;
    end else if (io_en) begin
      _T_44 <= _T_43;
    end
    if (reset) begin
      _T_45 <= 16'h0;
    end else if (io_en) begin
      _T_45 <= _T_44;
    end
    if (reset) begin
      _T_46 <= 16'h0;
    end else if (io_en) begin
      _T_46 <= _T_45;
    end
    if (reset) begin
      _T_47 <= 16'h0;
    end else if (io_en) begin
      _T_47 <= _T_46;
    end
    if (reset) begin
      _T_48 <= 16'h0;
    end else if (io_en) begin
      _T_48 <= _T_47;
    end
    if (reset) begin
      _T_49 <= 16'h0;
    end else if (io_en) begin
      _T_49 <= _T_48;
    end
    if (reset) begin
      _T_50 <= 16'h0;
    end else if (io_en) begin
      _T_50 <= _T_49;
    end
    if (reset) begin
      _T_51 <= 16'h0;
    end else if (io_en) begin
      _T_51 <= _T_50;
    end
    if (reset) begin
      _T_52 <= 16'h0;
    end else if (io_en) begin
      _T_52 <= _T_51;
    end
    if (reset) begin
      _T_53 <= 16'h0;
    end else if (io_en) begin
      _T_53 <= _T_52;
    end
    if (reset) begin
      _T_54 <= 16'h0;
    end else if (io_en) begin
      _T_54 <= _T_53;
    end
    if (reset) begin
      _T_55 <= 16'h0;
    end else if (io_en) begin
      _T_55 <= _T_54;
    end
    if (reset) begin
      _T_56 <= 16'h0;
    end else if (io_en) begin
      _T_56 <= _T_55;
    end
    if (reset) begin
      _T_57 <= 16'h0;
    end else if (io_en) begin
      _T_57 <= _T_56;
    end
    if (reset) begin
      _T_58 <= 16'h0;
    end else if (io_en) begin
      _T_58 <= _T_57;
    end
    if (reset) begin
      _T_59 <= 16'h0;
    end else if (io_en) begin
      _T_59 <= _T_58;
    end
    if (reset) begin
      _T_60 <= 16'h0;
    end else if (io_en) begin
      _T_60 <= _T_59;
    end
    if (reset) begin
      _T_61 <= 16'h0;
    end else if (io_en) begin
      _T_61 <= _T_60;
    end
    if (reset) begin
      _T_62 <= 16'h0;
    end else if (io_en) begin
      _T_62 <= _T_61;
    end
    if (reset) begin
      _T_63 <= 16'h0;
    end else if (io_en) begin
      _T_63 <= _T_62;
    end
    if (reset) begin
      _T_64 <= 16'h0;
    end else if (io_en) begin
      _T_64 <= _T_63;
    end
    if (reset) begin
      _T_65 <= 16'h0;
    end else if (io_en) begin
      _T_65 <= _T_64;
    end
    if (reset) begin
      _T_66 <= 16'h0;
    end else if (io_en) begin
      _T_66 <= _T_65;
    end
    if (reset) begin
      _T_67 <= 16'h0;
    end else if (io_en) begin
      _T_67 <= _T_66;
    end
    if (reset) begin
      _T_68 <= 16'h0;
    end else if (io_en) begin
      _T_68 <= _T_67;
    end
    if (reset) begin
      _T_69 <= 16'h0;
    end else if (io_en) begin
      _T_69 <= _T_68;
    end
    if (reset) begin
      _T_70 <= 16'h0;
    end else if (io_en) begin
      _T_70 <= _T_69;
    end
    if (reset) begin
      _T_71 <= 16'h0;
    end else if (io_en) begin
      _T_71 <= _T_70;
    end
    if (reset) begin
      _T_72 <= 16'h0;
    end else if (io_en) begin
      _T_72 <= _T_71;
    end
    if (reset) begin
      _T_73 <= 16'h0;
    end else if (io_en) begin
      _T_73 <= _T_72;
    end
    if (reset) begin
      _T_74 <= 16'h0;
    end else if (io_en) begin
      _T_74 <= _T_73;
    end
    if (reset) begin
      _T_75 <= 16'h0;
    end else if (io_en) begin
      _T_75 <= _T_74;
    end
    if (reset) begin
      _T_76 <= 16'h0;
    end else if (io_en) begin
      _T_76 <= _T_75;
    end
    if (reset) begin
      _T_77 <= 16'h0;
    end else if (io_en) begin
      _T_77 <= _T_76;
    end
    if (reset) begin
      _T_78 <= 16'h0;
    end else if (io_en) begin
      _T_78 <= _T_77;
    end
    if (reset) begin
      _T_79 <= 16'h0;
    end else if (io_en) begin
      _T_79 <= _T_78;
    end
    if (reset) begin
      _T_80 <= 16'h0;
    end else if (io_en) begin
      _T_80 <= _T_79;
    end
    if (reset) begin
      _T_81 <= 16'h0;
    end else if (io_en) begin
      _T_81 <= _T_80;
    end
    if (reset) begin
      _T_82 <= 16'h0;
    end else if (io_en) begin
      _T_82 <= _T_81;
    end
    if (reset) begin
      _T_83 <= 16'h0;
    end else if (io_en) begin
      _T_83 <= _T_82;
    end
    if (reset) begin
      _T_84 <= 16'h0;
    end else if (io_en) begin
      _T_84 <= _T_83;
    end
    if (reset) begin
      _T_85 <= 16'h0;
    end else if (io_en) begin
      _T_85 <= _T_84;
    end
    if (reset) begin
      _T_86 <= 16'h0;
    end else if (io_en) begin
      _T_86 <= _T_85;
    end
    if (reset) begin
      _T_87 <= 16'h0;
    end else if (io_en) begin
      _T_87 <= _T_86;
    end
    if (reset) begin
      _T_88 <= 16'h0;
    end else if (io_en) begin
      _T_88 <= _T_87;
    end
    if (reset) begin
      _T_89 <= 16'h0;
    end else if (io_en) begin
      _T_89 <= _T_88;
    end
    if (reset) begin
      _T_90 <= 16'h0;
    end else if (io_en) begin
      _T_90 <= _T_89;
    end
    if (reset) begin
      _T_91 <= 16'h0;
    end else if (io_en) begin
      _T_91 <= _T_90;
    end
    if (reset) begin
      _T_92 <= 16'h0;
    end else if (io_en) begin
      _T_92 <= _T_91;
    end
    if (reset) begin
      _T_93 <= 16'h0;
    end else if (io_en) begin
      _T_93 <= _T_92;
    end
    if (reset) begin
      _T_94 <= 16'h0;
    end else if (io_en) begin
      _T_94 <= _T_93;
    end
    if (reset) begin
      _T_95 <= 16'h0;
    end else if (io_en) begin
      _T_95 <= _T_94;
    end
    if (reset) begin
      _T_96 <= 16'h0;
    end else if (io_en) begin
      _T_96 <= _T_95;
    end
    if (reset) begin
      _T_97 <= 16'h0;
    end else if (io_en) begin
      _T_97 <= _T_96;
    end
    if (reset) begin
      _T_98 <= 16'h0;
    end else if (io_en) begin
      _T_98 <= _T_97;
    end
    if (reset) begin
      _T_99 <= 16'h0;
    end else if (io_en) begin
      _T_99 <= _T_98;
    end
    if (reset) begin
      _T_100 <= 16'h0;
    end else if (io_en) begin
      _T_100 <= _T_99;
    end
    if (reset) begin
      _T_101 <= 16'h0;
    end else if (io_en) begin
      _T_101 <= _T_100;
    end
    if (reset) begin
      _T_102 <= 16'h0;
    end else if (io_en) begin
      _T_102 <= _T_101;
    end
    if (reset) begin
      _T_103 <= 16'h0;
    end else if (io_en) begin
      _T_103 <= _T_102;
    end
    if (reset) begin
      _T_104 <= 16'h0;
    end else if (io_en) begin
      _T_104 <= _T_103;
    end
    if (reset) begin
      _T_105 <= 16'h0;
    end else if (io_en) begin
      _T_105 <= _T_104;
    end
    if (reset) begin
      _T_106 <= 16'h0;
    end else if (io_en) begin
      _T_106 <= _T_105;
    end
    if (reset) begin
      _T_107 <= 16'h0;
    end else if (io_en) begin
      _T_107 <= _T_106;
    end
    if (reset) begin
      _T_108 <= 16'h0;
    end else if (io_en) begin
      _T_108 <= _T_107;
    end
    if (reset) begin
      _T_109 <= 16'h0;
    end else if (io_en) begin
      _T_109 <= _T_108;
    end
    if (reset) begin
      _T_110 <= 16'h0;
    end else if (io_en) begin
      _T_110 <= _T_109;
    end
    if (reset) begin
      _T_111 <= 16'h0;
    end else if (io_en) begin
      _T_111 <= _T_110;
    end
    if (reset) begin
      _T_112 <= 16'h0;
    end else if (io_en) begin
      _T_112 <= _T_111;
    end
    if (reset) begin
      _T_113 <= 16'h0;
    end else if (io_en) begin
      _T_113 <= _T_112;
    end
    if (reset) begin
      _T_114 <= 16'h0;
    end else if (io_en) begin
      _T_114 <= _T_113;
    end
    if (reset) begin
      _T_115 <= 16'h0;
    end else if (io_en) begin
      _T_115 <= _T_114;
    end
    if (reset) begin
      _T_116 <= 16'h0;
    end else if (io_en) begin
      _T_116 <= _T_115;
    end
    if (reset) begin
      _T_117 <= 16'h0;
    end else if (io_en) begin
      _T_117 <= _T_116;
    end
    if (reset) begin
      _T_118 <= 16'h0;
    end else if (io_en) begin
      _T_118 <= _T_117;
    end
    if (reset) begin
      _T_119 <= 16'h0;
    end else if (io_en) begin
      _T_119 <= _T_118;
    end
  end
endmodule
module Mac_103(
  input           clock,
  input           reset,
  input  [1919:0] io_a,
  input  [1919:0] io_b,
  input           io_rdy,
  output [31:0]   io_q,
  output          io_v
);
  wire [15:0] a_0;
  wire [15:0] b_0;
  wire [15:0] a_1;
  wire [15:0] b_1;
  wire [15:0] a_2;
  wire [15:0] b_2;
  wire [15:0] a_3;
  wire [15:0] b_3;
  wire [15:0] a_4;
  wire [15:0] b_4;
  wire [15:0] a_5;
  wire [15:0] b_5;
  wire [15:0] a_6;
  wire [15:0] b_6;
  wire [15:0] a_7;
  wire [15:0] b_7;
  wire [15:0] a_8;
  wire [15:0] b_8;
  wire [15:0] a_9;
  wire [15:0] b_9;
  wire [15:0] a_10;
  wire [15:0] b_10;
  wire [15:0] a_11;
  wire [15:0] b_11;
  wire [15:0] a_12;
  wire [15:0] b_12;
  wire [15:0] a_13;
  wire [15:0] b_13;
  wire [15:0] a_14;
  wire [15:0] b_14;
  wire [15:0] a_15;
  wire [15:0] b_15;
  wire [15:0] a_16;
  wire [15:0] b_16;
  wire [15:0] a_17;
  wire [15:0] b_17;
  wire [15:0] a_18;
  wire [15:0] b_18;
  wire [15:0] a_19;
  wire [15:0] b_19;
  wire [15:0] a_20;
  wire [15:0] b_20;
  wire [15:0] a_21;
  wire [15:0] b_21;
  wire [15:0] a_22;
  wire [15:0] b_22;
  wire [15:0] a_23;
  wire [15:0] b_23;
  wire [15:0] a_24;
  wire [15:0] b_24;
  wire [15:0] a_25;
  wire [15:0] b_25;
  wire [15:0] a_26;
  wire [15:0] b_26;
  wire [15:0] a_27;
  wire [15:0] b_27;
  wire [15:0] a_28;
  wire [15:0] b_28;
  wire [15:0] a_29;
  wire [15:0] b_29;
  wire [15:0] a_30;
  wire [15:0] b_30;
  wire [15:0] a_31;
  wire [15:0] b_31;
  wire [15:0] a_32;
  wire [15:0] b_32;
  wire [15:0] a_33;
  wire [15:0] b_33;
  wire [15:0] a_34;
  wire [15:0] b_34;
  wire [15:0] a_35;
  wire [15:0] b_35;
  wire [15:0] a_36;
  wire [15:0] b_36;
  wire [15:0] a_37;
  wire [15:0] b_37;
  wire [15:0] a_38;
  wire [15:0] b_38;
  wire [15:0] a_39;
  wire [15:0] b_39;
  wire [15:0] a_40;
  wire [15:0] b_40;
  wire [15:0] a_41;
  wire [15:0] b_41;
  wire [15:0] a_42;
  wire [15:0] b_42;
  wire [15:0] a_43;
  wire [15:0] b_43;
  wire [15:0] a_44;
  wire [15:0] b_44;
  wire [15:0] a_45;
  wire [15:0] b_45;
  wire [15:0] a_46;
  wire [15:0] b_46;
  wire [15:0] a_47;
  wire [15:0] b_47;
  wire [15:0] a_48;
  wire [15:0] b_48;
  wire [15:0] a_49;
  wire [15:0] b_49;
  wire [15:0] a_50;
  wire [15:0] b_50;
  wire [15:0] a_51;
  wire [15:0] b_51;
  wire [15:0] a_52;
  wire [15:0] b_52;
  wire [15:0] a_53;
  wire [15:0] b_53;
  wire [15:0] a_54;
  wire [15:0] b_54;
  wire [15:0] a_55;
  wire [15:0] b_55;
  wire [15:0] a_56;
  wire [15:0] b_56;
  wire [15:0] a_57;
  wire [15:0] b_57;
  wire [15:0] a_58;
  wire [15:0] b_58;
  wire [15:0] a_59;
  wire [15:0] b_59;
  wire [15:0] a_60;
  wire [15:0] b_60;
  wire [15:0] a_61;
  wire [15:0] b_61;
  wire [15:0] a_62;
  wire [15:0] b_62;
  wire [15:0] a_63;
  wire [15:0] b_63;
  wire [15:0] a_64;
  wire [15:0] b_64;
  wire [15:0] a_65;
  wire [15:0] b_65;
  wire [15:0] a_66;
  wire [15:0] b_66;
  wire [15:0] a_67;
  wire [15:0] b_67;
  wire [15:0] a_68;
  wire [15:0] b_68;
  wire [15:0] a_69;
  wire [15:0] b_69;
  wire [15:0] a_70;
  wire [15:0] b_70;
  wire [15:0] a_71;
  wire [15:0] b_71;
  wire [15:0] a_72;
  wire [15:0] b_72;
  wire [15:0] a_73;
  wire [15:0] b_73;
  wire [15:0] a_74;
  wire [15:0] b_74;
  wire [15:0] a_75;
  wire [15:0] b_75;
  wire [15:0] a_76;
  wire [15:0] b_76;
  wire [15:0] a_77;
  wire [15:0] b_77;
  wire [15:0] a_78;
  wire [15:0] b_78;
  wire [15:0] a_79;
  wire [15:0] b_79;
  wire [15:0] a_80;
  wire [15:0] b_80;
  wire [15:0] a_81;
  wire [15:0] b_81;
  wire [15:0] a_82;
  wire [15:0] b_82;
  wire [15:0] a_83;
  wire [15:0] b_83;
  wire [15:0] a_84;
  wire [15:0] b_84;
  wire [15:0] a_85;
  wire [15:0] b_85;
  wire [15:0] a_86;
  wire [15:0] b_86;
  wire [15:0] a_87;
  wire [15:0] b_87;
  wire [15:0] a_88;
  wire [15:0] b_88;
  wire [15:0] a_89;
  wire [15:0] b_89;
  wire [15:0] a_90;
  wire [15:0] b_90;
  wire [15:0] a_91;
  wire [15:0] b_91;
  wire [15:0] a_92;
  wire [15:0] b_92;
  wire [15:0] a_93;
  wire [15:0] b_93;
  wire [15:0] a_94;
  wire [15:0] b_94;
  wire [15:0] a_95;
  wire [15:0] b_95;
  wire [15:0] a_96;
  wire [15:0] b_96;
  wire [15:0] a_97;
  wire [15:0] b_97;
  wire [15:0] a_98;
  wire [15:0] b_98;
  wire [15:0] a_99;
  wire [15:0] b_99;
  wire [15:0] a_100;
  wire [15:0] b_100;
  wire [15:0] a_101;
  wire [15:0] b_101;
  wire [15:0] a_102;
  wire [15:0] b_102;
  wire [15:0] a_103;
  wire [15:0] b_103;
  wire [15:0] a_104;
  wire [15:0] b_104;
  wire [15:0] a_105;
  wire [15:0] b_105;
  wire [15:0] a_106;
  wire [15:0] b_106;
  wire [15:0] a_107;
  wire [15:0] b_107;
  wire [15:0] a_108;
  wire [15:0] b_108;
  wire [15:0] a_109;
  wire [15:0] b_109;
  wire [15:0] a_110;
  wire [15:0] b_110;
  wire [15:0] a_111;
  wire [15:0] b_111;
  wire [15:0] a_112;
  wire [15:0] b_112;
  wire [15:0] a_113;
  wire [15:0] b_113;
  wire [15:0] a_114;
  wire [15:0] b_114;
  wire [15:0] a_115;
  wire [15:0] b_115;
  wire [15:0] a_116;
  wire [15:0] b_116;
  wire [15:0] a_117;
  wire [15:0] b_117;
  wire [15:0] a_118;
  wire [15:0] b_118;
  wire [15:0] a_119;
  wire [15:0] b_119;
  reg [31:0] sum;
  reg [31:0] _RAND_0;
  reg [6:0] i;
  reg [31:0] _RAND_1;
  wire  _T_243;
  wire  _T_244;
  wire [15:0] _GEN_1;
  wire [15:0] _GEN_2;
  wire [15:0] _GEN_3;
  wire [15:0] _GEN_4;
  wire [15:0] _GEN_5;
  wire [15:0] _GEN_6;
  wire [15:0] _GEN_7;
  wire [15:0] _GEN_8;
  wire [15:0] _GEN_9;
  wire [15:0] _GEN_10;
  wire [15:0] _GEN_11;
  wire [15:0] _GEN_12;
  wire [15:0] _GEN_13;
  wire [15:0] _GEN_14;
  wire [15:0] _GEN_15;
  wire [15:0] _GEN_16;
  wire [15:0] _GEN_17;
  wire [15:0] _GEN_18;
  wire [15:0] _GEN_19;
  wire [15:0] _GEN_20;
  wire [15:0] _GEN_21;
  wire [15:0] _GEN_22;
  wire [15:0] _GEN_23;
  wire [15:0] _GEN_24;
  wire [15:0] _GEN_25;
  wire [15:0] _GEN_26;
  wire [15:0] _GEN_27;
  wire [15:0] _GEN_28;
  wire [15:0] _GEN_29;
  wire [15:0] _GEN_30;
  wire [15:0] _GEN_31;
  wire [15:0] _GEN_32;
  wire [15:0] _GEN_33;
  wire [15:0] _GEN_34;
  wire [15:0] _GEN_35;
  wire [15:0] _GEN_36;
  wire [15:0] _GEN_37;
  wire [15:0] _GEN_38;
  wire [15:0] _GEN_39;
  wire [15:0] _GEN_40;
  wire [15:0] _GEN_41;
  wire [15:0] _GEN_42;
  wire [15:0] _GEN_43;
  wire [15:0] _GEN_44;
  wire [15:0] _GEN_45;
  wire [15:0] _GEN_46;
  wire [15:0] _GEN_47;
  wire [15:0] _GEN_48;
  wire [15:0] _GEN_49;
  wire [15:0] _GEN_50;
  wire [15:0] _GEN_51;
  wire [15:0] _GEN_52;
  wire [15:0] _GEN_53;
  wire [15:0] _GEN_54;
  wire [15:0] _GEN_55;
  wire [15:0] _GEN_56;
  wire [15:0] _GEN_57;
  wire [15:0] _GEN_58;
  wire [15:0] _GEN_59;
  wire [15:0] _GEN_60;
  wire [15:0] _GEN_61;
  wire [15:0] _GEN_62;
  wire [15:0] _GEN_63;
  wire [15:0] _GEN_64;
  wire [15:0] _GEN_65;
  wire [15:0] _GEN_66;
  wire [15:0] _GEN_67;
  wire [15:0] _GEN_68;
  wire [15:0] _GEN_69;
  wire [15:0] _GEN_70;
  wire [15:0] _GEN_71;
  wire [15:0] _GEN_72;
  wire [15:0] _GEN_73;
  wire [15:0] _GEN_74;
  wire [15:0] _GEN_75;
  wire [15:0] _GEN_76;
  wire [15:0] _GEN_77;
  wire [15:0] _GEN_78;
  wire [15:0] _GEN_79;
  wire [15:0] _GEN_80;
  wire [15:0] _GEN_81;
  wire [15:0] _GEN_82;
  wire [15:0] _GEN_83;
  wire [15:0] _GEN_84;
  wire [15:0] _GEN_85;
  wire [15:0] _GEN_86;
  wire [15:0] _GEN_87;
  wire [15:0] _GEN_88;
  wire [15:0] _GEN_89;
  wire [15:0] _GEN_90;
  wire [15:0] _GEN_91;
  wire [15:0] _GEN_92;
  wire [15:0] _GEN_93;
  wire [15:0] _GEN_94;
  wire [15:0] _GEN_95;
  wire [15:0] _GEN_96;
  wire [15:0] _GEN_97;
  wire [15:0] _GEN_98;
  wire [15:0] _GEN_99;
  wire [15:0] _GEN_100;
  wire [15:0] _GEN_101;
  wire [15:0] _GEN_102;
  wire [15:0] _GEN_103;
  wire [15:0] _GEN_104;
  wire [15:0] _GEN_105;
  wire [15:0] _GEN_106;
  wire [15:0] _GEN_107;
  wire [15:0] _GEN_108;
  wire [15:0] _GEN_109;
  wire [15:0] _GEN_110;
  wire [15:0] _GEN_111;
  wire [15:0] _GEN_112;
  wire [15:0] _GEN_113;
  wire [15:0] _GEN_114;
  wire [15:0] _GEN_115;
  wire [15:0] _GEN_116;
  wire [15:0] _GEN_117;
  wire [15:0] _GEN_118;
  wire [15:0] _GEN_119;
  wire [15:0] _GEN_121;
  wire [15:0] _GEN_122;
  wire [15:0] _GEN_123;
  wire [15:0] _GEN_124;
  wire [15:0] _GEN_125;
  wire [15:0] _GEN_126;
  wire [15:0] _GEN_127;
  wire [15:0] _GEN_128;
  wire [15:0] _GEN_129;
  wire [15:0] _GEN_130;
  wire [15:0] _GEN_131;
  wire [15:0] _GEN_132;
  wire [15:0] _GEN_133;
  wire [15:0] _GEN_134;
  wire [15:0] _GEN_135;
  wire [15:0] _GEN_136;
  wire [15:0] _GEN_137;
  wire [15:0] _GEN_138;
  wire [15:0] _GEN_139;
  wire [15:0] _GEN_140;
  wire [15:0] _GEN_141;
  wire [15:0] _GEN_142;
  wire [15:0] _GEN_143;
  wire [15:0] _GEN_144;
  wire [15:0] _GEN_145;
  wire [15:0] _GEN_146;
  wire [15:0] _GEN_147;
  wire [15:0] _GEN_148;
  wire [15:0] _GEN_149;
  wire [15:0] _GEN_150;
  wire [15:0] _GEN_151;
  wire [15:0] _GEN_152;
  wire [15:0] _GEN_153;
  wire [15:0] _GEN_154;
  wire [15:0] _GEN_155;
  wire [15:0] _GEN_156;
  wire [15:0] _GEN_157;
  wire [15:0] _GEN_158;
  wire [15:0] _GEN_159;
  wire [15:0] _GEN_160;
  wire [15:0] _GEN_161;
  wire [15:0] _GEN_162;
  wire [15:0] _GEN_163;
  wire [15:0] _GEN_164;
  wire [15:0] _GEN_165;
  wire [15:0] _GEN_166;
  wire [15:0] _GEN_167;
  wire [15:0] _GEN_168;
  wire [15:0] _GEN_169;
  wire [15:0] _GEN_170;
  wire [15:0] _GEN_171;
  wire [15:0] _GEN_172;
  wire [15:0] _GEN_173;
  wire [15:0] _GEN_174;
  wire [15:0] _GEN_175;
  wire [15:0] _GEN_176;
  wire [15:0] _GEN_177;
  wire [15:0] _GEN_178;
  wire [15:0] _GEN_179;
  wire [15:0] _GEN_180;
  wire [15:0] _GEN_181;
  wire [15:0] _GEN_182;
  wire [15:0] _GEN_183;
  wire [15:0] _GEN_184;
  wire [15:0] _GEN_185;
  wire [15:0] _GEN_186;
  wire [15:0] _GEN_187;
  wire [15:0] _GEN_188;
  wire [15:0] _GEN_189;
  wire [15:0] _GEN_190;
  wire [15:0] _GEN_191;
  wire [15:0] _GEN_192;
  wire [15:0] _GEN_193;
  wire [15:0] _GEN_194;
  wire [15:0] _GEN_195;
  wire [15:0] _GEN_196;
  wire [15:0] _GEN_197;
  wire [15:0] _GEN_198;
  wire [15:0] _GEN_199;
  wire [15:0] _GEN_200;
  wire [15:0] _GEN_201;
  wire [15:0] _GEN_202;
  wire [15:0] _GEN_203;
  wire [15:0] _GEN_204;
  wire [15:0] _GEN_205;
  wire [15:0] _GEN_206;
  wire [15:0] _GEN_207;
  wire [15:0] _GEN_208;
  wire [15:0] _GEN_209;
  wire [15:0] _GEN_210;
  wire [15:0] _GEN_211;
  wire [15:0] _GEN_212;
  wire [15:0] _GEN_213;
  wire [15:0] _GEN_214;
  wire [15:0] _GEN_215;
  wire [15:0] _GEN_216;
  wire [15:0] _GEN_217;
  wire [15:0] _GEN_218;
  wire [15:0] _GEN_219;
  wire [15:0] _GEN_220;
  wire [15:0] _GEN_221;
  wire [15:0] _GEN_222;
  wire [15:0] _GEN_223;
  wire [15:0] _GEN_224;
  wire [15:0] _GEN_225;
  wire [15:0] _GEN_226;
  wire [15:0] _GEN_227;
  wire [15:0] _GEN_228;
  wire [15:0] _GEN_229;
  wire [15:0] _GEN_230;
  wire [15:0] _GEN_231;
  wire [15:0] _GEN_232;
  wire [15:0] _GEN_233;
  wire [15:0] _GEN_234;
  wire [15:0] _GEN_235;
  wire [15:0] _GEN_236;
  wire [15:0] _GEN_237;
  wire [15:0] _GEN_238;
  wire [15:0] _GEN_239;
  wire [31:0] _T_240;
  wire [32:0] _T_241;
  wire [7:0] _T_242;
  wire [7:0] _GEN_240;
  wire [32:0] _GEN_241;
  wire [7:0] _GEN_242;
  wire [31:0] _GEN_244;
  wire [32:0] _GEN_245;
  wire [32:0] _GEN_246;
  wire [7:0] _GEN_247;
  assign a_0 = io_a[15:0];
  assign b_0 = io_b[15:0];
  assign a_1 = io_a[31:16];
  assign b_1 = io_b[31:16];
  assign a_2 = io_a[47:32];
  assign b_2 = io_b[47:32];
  assign a_3 = io_a[63:48];
  assign b_3 = io_b[63:48];
  assign a_4 = io_a[79:64];
  assign b_4 = io_b[79:64];
  assign a_5 = io_a[95:80];
  assign b_5 = io_b[95:80];
  assign a_6 = io_a[111:96];
  assign b_6 = io_b[111:96];
  assign a_7 = io_a[127:112];
  assign b_7 = io_b[127:112];
  assign a_8 = io_a[143:128];
  assign b_8 = io_b[143:128];
  assign a_9 = io_a[159:144];
  assign b_9 = io_b[159:144];
  assign a_10 = io_a[175:160];
  assign b_10 = io_b[175:160];
  assign a_11 = io_a[191:176];
  assign b_11 = io_b[191:176];
  assign a_12 = io_a[207:192];
  assign b_12 = io_b[207:192];
  assign a_13 = io_a[223:208];
  assign b_13 = io_b[223:208];
  assign a_14 = io_a[239:224];
  assign b_14 = io_b[239:224];
  assign a_15 = io_a[255:240];
  assign b_15 = io_b[255:240];
  assign a_16 = io_a[271:256];
  assign b_16 = io_b[271:256];
  assign a_17 = io_a[287:272];
  assign b_17 = io_b[287:272];
  assign a_18 = io_a[303:288];
  assign b_18 = io_b[303:288];
  assign a_19 = io_a[319:304];
  assign b_19 = io_b[319:304];
  assign a_20 = io_a[335:320];
  assign b_20 = io_b[335:320];
  assign a_21 = io_a[351:336];
  assign b_21 = io_b[351:336];
  assign a_22 = io_a[367:352];
  assign b_22 = io_b[367:352];
  assign a_23 = io_a[383:368];
  assign b_23 = io_b[383:368];
  assign a_24 = io_a[399:384];
  assign b_24 = io_b[399:384];
  assign a_25 = io_a[415:400];
  assign b_25 = io_b[415:400];
  assign a_26 = io_a[431:416];
  assign b_26 = io_b[431:416];
  assign a_27 = io_a[447:432];
  assign b_27 = io_b[447:432];
  assign a_28 = io_a[463:448];
  assign b_28 = io_b[463:448];
  assign a_29 = io_a[479:464];
  assign b_29 = io_b[479:464];
  assign a_30 = io_a[495:480];
  assign b_30 = io_b[495:480];
  assign a_31 = io_a[511:496];
  assign b_31 = io_b[511:496];
  assign a_32 = io_a[527:512];
  assign b_32 = io_b[527:512];
  assign a_33 = io_a[543:528];
  assign b_33 = io_b[543:528];
  assign a_34 = io_a[559:544];
  assign b_34 = io_b[559:544];
  assign a_35 = io_a[575:560];
  assign b_35 = io_b[575:560];
  assign a_36 = io_a[591:576];
  assign b_36 = io_b[591:576];
  assign a_37 = io_a[607:592];
  assign b_37 = io_b[607:592];
  assign a_38 = io_a[623:608];
  assign b_38 = io_b[623:608];
  assign a_39 = io_a[639:624];
  assign b_39 = io_b[639:624];
  assign a_40 = io_a[655:640];
  assign b_40 = io_b[655:640];
  assign a_41 = io_a[671:656];
  assign b_41 = io_b[671:656];
  assign a_42 = io_a[687:672];
  assign b_42 = io_b[687:672];
  assign a_43 = io_a[703:688];
  assign b_43 = io_b[703:688];
  assign a_44 = io_a[719:704];
  assign b_44 = io_b[719:704];
  assign a_45 = io_a[735:720];
  assign b_45 = io_b[735:720];
  assign a_46 = io_a[751:736];
  assign b_46 = io_b[751:736];
  assign a_47 = io_a[767:752];
  assign b_47 = io_b[767:752];
  assign a_48 = io_a[783:768];
  assign b_48 = io_b[783:768];
  assign a_49 = io_a[799:784];
  assign b_49 = io_b[799:784];
  assign a_50 = io_a[815:800];
  assign b_50 = io_b[815:800];
  assign a_51 = io_a[831:816];
  assign b_51 = io_b[831:816];
  assign a_52 = io_a[847:832];
  assign b_52 = io_b[847:832];
  assign a_53 = io_a[863:848];
  assign b_53 = io_b[863:848];
  assign a_54 = io_a[879:864];
  assign b_54 = io_b[879:864];
  assign a_55 = io_a[895:880];
  assign b_55 = io_b[895:880];
  assign a_56 = io_a[911:896];
  assign b_56 = io_b[911:896];
  assign a_57 = io_a[927:912];
  assign b_57 = io_b[927:912];
  assign a_58 = io_a[943:928];
  assign b_58 = io_b[943:928];
  assign a_59 = io_a[959:944];
  assign b_59 = io_b[959:944];
  assign a_60 = io_a[975:960];
  assign b_60 = io_b[975:960];
  assign a_61 = io_a[991:976];
  assign b_61 = io_b[991:976];
  assign a_62 = io_a[1007:992];
  assign b_62 = io_b[1007:992];
  assign a_63 = io_a[1023:1008];
  assign b_63 = io_b[1023:1008];
  assign a_64 = io_a[1039:1024];
  assign b_64 = io_b[1039:1024];
  assign a_65 = io_a[1055:1040];
  assign b_65 = io_b[1055:1040];
  assign a_66 = io_a[1071:1056];
  assign b_66 = io_b[1071:1056];
  assign a_67 = io_a[1087:1072];
  assign b_67 = io_b[1087:1072];
  assign a_68 = io_a[1103:1088];
  assign b_68 = io_b[1103:1088];
  assign a_69 = io_a[1119:1104];
  assign b_69 = io_b[1119:1104];
  assign a_70 = io_a[1135:1120];
  assign b_70 = io_b[1135:1120];
  assign a_71 = io_a[1151:1136];
  assign b_71 = io_b[1151:1136];
  assign a_72 = io_a[1167:1152];
  assign b_72 = io_b[1167:1152];
  assign a_73 = io_a[1183:1168];
  assign b_73 = io_b[1183:1168];
  assign a_74 = io_a[1199:1184];
  assign b_74 = io_b[1199:1184];
  assign a_75 = io_a[1215:1200];
  assign b_75 = io_b[1215:1200];
  assign a_76 = io_a[1231:1216];
  assign b_76 = io_b[1231:1216];
  assign a_77 = io_a[1247:1232];
  assign b_77 = io_b[1247:1232];
  assign a_78 = io_a[1263:1248];
  assign b_78 = io_b[1263:1248];
  assign a_79 = io_a[1279:1264];
  assign b_79 = io_b[1279:1264];
  assign a_80 = io_a[1295:1280];
  assign b_80 = io_b[1295:1280];
  assign a_81 = io_a[1311:1296];
  assign b_81 = io_b[1311:1296];
  assign a_82 = io_a[1327:1312];
  assign b_82 = io_b[1327:1312];
  assign a_83 = io_a[1343:1328];
  assign b_83 = io_b[1343:1328];
  assign a_84 = io_a[1359:1344];
  assign b_84 = io_b[1359:1344];
  assign a_85 = io_a[1375:1360];
  assign b_85 = io_b[1375:1360];
  assign a_86 = io_a[1391:1376];
  assign b_86 = io_b[1391:1376];
  assign a_87 = io_a[1407:1392];
  assign b_87 = io_b[1407:1392];
  assign a_88 = io_a[1423:1408];
  assign b_88 = io_b[1423:1408];
  assign a_89 = io_a[1439:1424];
  assign b_89 = io_b[1439:1424];
  assign a_90 = io_a[1455:1440];
  assign b_90 = io_b[1455:1440];
  assign a_91 = io_a[1471:1456];
  assign b_91 = io_b[1471:1456];
  assign a_92 = io_a[1487:1472];
  assign b_92 = io_b[1487:1472];
  assign a_93 = io_a[1503:1488];
  assign b_93 = io_b[1503:1488];
  assign a_94 = io_a[1519:1504];
  assign b_94 = io_b[1519:1504];
  assign a_95 = io_a[1535:1520];
  assign b_95 = io_b[1535:1520];
  assign a_96 = io_a[1551:1536];
  assign b_96 = io_b[1551:1536];
  assign a_97 = io_a[1567:1552];
  assign b_97 = io_b[1567:1552];
  assign a_98 = io_a[1583:1568];
  assign b_98 = io_b[1583:1568];
  assign a_99 = io_a[1599:1584];
  assign b_99 = io_b[1599:1584];
  assign a_100 = io_a[1615:1600];
  assign b_100 = io_b[1615:1600];
  assign a_101 = io_a[1631:1616];
  assign b_101 = io_b[1631:1616];
  assign a_102 = io_a[1647:1632];
  assign b_102 = io_b[1647:1632];
  assign a_103 = io_a[1663:1648];
  assign b_103 = io_b[1663:1648];
  assign a_104 = io_a[1679:1664];
  assign b_104 = io_b[1679:1664];
  assign a_105 = io_a[1695:1680];
  assign b_105 = io_b[1695:1680];
  assign a_106 = io_a[1711:1696];
  assign b_106 = io_b[1711:1696];
  assign a_107 = io_a[1727:1712];
  assign b_107 = io_b[1727:1712];
  assign a_108 = io_a[1743:1728];
  assign b_108 = io_b[1743:1728];
  assign a_109 = io_a[1759:1744];
  assign b_109 = io_b[1759:1744];
  assign a_110 = io_a[1775:1760];
  assign b_110 = io_b[1775:1760];
  assign a_111 = io_a[1791:1776];
  assign b_111 = io_b[1791:1776];
  assign a_112 = io_a[1807:1792];
  assign b_112 = io_b[1807:1792];
  assign a_113 = io_a[1823:1808];
  assign b_113 = io_b[1823:1808];
  assign a_114 = io_a[1839:1824];
  assign b_114 = io_b[1839:1824];
  assign a_115 = io_a[1855:1840];
  assign b_115 = io_b[1855:1840];
  assign a_116 = io_a[1871:1856];
  assign b_116 = io_b[1871:1856];
  assign a_117 = io_a[1887:1872];
  assign b_117 = io_b[1887:1872];
  assign a_118 = io_a[1903:1888];
  assign b_118 = io_b[1903:1888];
  assign a_119 = io_a[1919:1904];
  assign b_119 = io_b[1919:1904];
  assign _T_243 = i == 7'h78;
  assign _T_244 = i != 7'h0;
  assign _GEN_1 = 7'h1 == i ? a_1 : a_0;
  assign _GEN_2 = 7'h2 == i ? a_2 : _GEN_1;
  assign _GEN_3 = 7'h3 == i ? a_3 : _GEN_2;
  assign _GEN_4 = 7'h4 == i ? a_4 : _GEN_3;
  assign _GEN_5 = 7'h5 == i ? a_5 : _GEN_4;
  assign _GEN_6 = 7'h6 == i ? a_6 : _GEN_5;
  assign _GEN_7 = 7'h7 == i ? a_7 : _GEN_6;
  assign _GEN_8 = 7'h8 == i ? a_8 : _GEN_7;
  assign _GEN_9 = 7'h9 == i ? a_9 : _GEN_8;
  assign _GEN_10 = 7'ha == i ? a_10 : _GEN_9;
  assign _GEN_11 = 7'hb == i ? a_11 : _GEN_10;
  assign _GEN_12 = 7'hc == i ? a_12 : _GEN_11;
  assign _GEN_13 = 7'hd == i ? a_13 : _GEN_12;
  assign _GEN_14 = 7'he == i ? a_14 : _GEN_13;
  assign _GEN_15 = 7'hf == i ? a_15 : _GEN_14;
  assign _GEN_16 = 7'h10 == i ? a_16 : _GEN_15;
  assign _GEN_17 = 7'h11 == i ? a_17 : _GEN_16;
  assign _GEN_18 = 7'h12 == i ? a_18 : _GEN_17;
  assign _GEN_19 = 7'h13 == i ? a_19 : _GEN_18;
  assign _GEN_20 = 7'h14 == i ? a_20 : _GEN_19;
  assign _GEN_21 = 7'h15 == i ? a_21 : _GEN_20;
  assign _GEN_22 = 7'h16 == i ? a_22 : _GEN_21;
  assign _GEN_23 = 7'h17 == i ? a_23 : _GEN_22;
  assign _GEN_24 = 7'h18 == i ? a_24 : _GEN_23;
  assign _GEN_25 = 7'h19 == i ? a_25 : _GEN_24;
  assign _GEN_26 = 7'h1a == i ? a_26 : _GEN_25;
  assign _GEN_27 = 7'h1b == i ? a_27 : _GEN_26;
  assign _GEN_28 = 7'h1c == i ? a_28 : _GEN_27;
  assign _GEN_29 = 7'h1d == i ? a_29 : _GEN_28;
  assign _GEN_30 = 7'h1e == i ? a_30 : _GEN_29;
  assign _GEN_31 = 7'h1f == i ? a_31 : _GEN_30;
  assign _GEN_32 = 7'h20 == i ? a_32 : _GEN_31;
  assign _GEN_33 = 7'h21 == i ? a_33 : _GEN_32;
  assign _GEN_34 = 7'h22 == i ? a_34 : _GEN_33;
  assign _GEN_35 = 7'h23 == i ? a_35 : _GEN_34;
  assign _GEN_36 = 7'h24 == i ? a_36 : _GEN_35;
  assign _GEN_37 = 7'h25 == i ? a_37 : _GEN_36;
  assign _GEN_38 = 7'h26 == i ? a_38 : _GEN_37;
  assign _GEN_39 = 7'h27 == i ? a_39 : _GEN_38;
  assign _GEN_40 = 7'h28 == i ? a_40 : _GEN_39;
  assign _GEN_41 = 7'h29 == i ? a_41 : _GEN_40;
  assign _GEN_42 = 7'h2a == i ? a_42 : _GEN_41;
  assign _GEN_43 = 7'h2b == i ? a_43 : _GEN_42;
  assign _GEN_44 = 7'h2c == i ? a_44 : _GEN_43;
  assign _GEN_45 = 7'h2d == i ? a_45 : _GEN_44;
  assign _GEN_46 = 7'h2e == i ? a_46 : _GEN_45;
  assign _GEN_47 = 7'h2f == i ? a_47 : _GEN_46;
  assign _GEN_48 = 7'h30 == i ? a_48 : _GEN_47;
  assign _GEN_49 = 7'h31 == i ? a_49 : _GEN_48;
  assign _GEN_50 = 7'h32 == i ? a_50 : _GEN_49;
  assign _GEN_51 = 7'h33 == i ? a_51 : _GEN_50;
  assign _GEN_52 = 7'h34 == i ? a_52 : _GEN_51;
  assign _GEN_53 = 7'h35 == i ? a_53 : _GEN_52;
  assign _GEN_54 = 7'h36 == i ? a_54 : _GEN_53;
  assign _GEN_55 = 7'h37 == i ? a_55 : _GEN_54;
  assign _GEN_56 = 7'h38 == i ? a_56 : _GEN_55;
  assign _GEN_57 = 7'h39 == i ? a_57 : _GEN_56;
  assign _GEN_58 = 7'h3a == i ? a_58 : _GEN_57;
  assign _GEN_59 = 7'h3b == i ? a_59 : _GEN_58;
  assign _GEN_60 = 7'h3c == i ? a_60 : _GEN_59;
  assign _GEN_61 = 7'h3d == i ? a_61 : _GEN_60;
  assign _GEN_62 = 7'h3e == i ? a_62 : _GEN_61;
  assign _GEN_63 = 7'h3f == i ? a_63 : _GEN_62;
  assign _GEN_64 = 7'h40 == i ? a_64 : _GEN_63;
  assign _GEN_65 = 7'h41 == i ? a_65 : _GEN_64;
  assign _GEN_66 = 7'h42 == i ? a_66 : _GEN_65;
  assign _GEN_67 = 7'h43 == i ? a_67 : _GEN_66;
  assign _GEN_68 = 7'h44 == i ? a_68 : _GEN_67;
  assign _GEN_69 = 7'h45 == i ? a_69 : _GEN_68;
  assign _GEN_70 = 7'h46 == i ? a_70 : _GEN_69;
  assign _GEN_71 = 7'h47 == i ? a_71 : _GEN_70;
  assign _GEN_72 = 7'h48 == i ? a_72 : _GEN_71;
  assign _GEN_73 = 7'h49 == i ? a_73 : _GEN_72;
  assign _GEN_74 = 7'h4a == i ? a_74 : _GEN_73;
  assign _GEN_75 = 7'h4b == i ? a_75 : _GEN_74;
  assign _GEN_76 = 7'h4c == i ? a_76 : _GEN_75;
  assign _GEN_77 = 7'h4d == i ? a_77 : _GEN_76;
  assign _GEN_78 = 7'h4e == i ? a_78 : _GEN_77;
  assign _GEN_79 = 7'h4f == i ? a_79 : _GEN_78;
  assign _GEN_80 = 7'h50 == i ? a_80 : _GEN_79;
  assign _GEN_81 = 7'h51 == i ? a_81 : _GEN_80;
  assign _GEN_82 = 7'h52 == i ? a_82 : _GEN_81;
  assign _GEN_83 = 7'h53 == i ? a_83 : _GEN_82;
  assign _GEN_84 = 7'h54 == i ? a_84 : _GEN_83;
  assign _GEN_85 = 7'h55 == i ? a_85 : _GEN_84;
  assign _GEN_86 = 7'h56 == i ? a_86 : _GEN_85;
  assign _GEN_87 = 7'h57 == i ? a_87 : _GEN_86;
  assign _GEN_88 = 7'h58 == i ? a_88 : _GEN_87;
  assign _GEN_89 = 7'h59 == i ? a_89 : _GEN_88;
  assign _GEN_90 = 7'h5a == i ? a_90 : _GEN_89;
  assign _GEN_91 = 7'h5b == i ? a_91 : _GEN_90;
  assign _GEN_92 = 7'h5c == i ? a_92 : _GEN_91;
  assign _GEN_93 = 7'h5d == i ? a_93 : _GEN_92;
  assign _GEN_94 = 7'h5e == i ? a_94 : _GEN_93;
  assign _GEN_95 = 7'h5f == i ? a_95 : _GEN_94;
  assign _GEN_96 = 7'h60 == i ? a_96 : _GEN_95;
  assign _GEN_97 = 7'h61 == i ? a_97 : _GEN_96;
  assign _GEN_98 = 7'h62 == i ? a_98 : _GEN_97;
  assign _GEN_99 = 7'h63 == i ? a_99 : _GEN_98;
  assign _GEN_100 = 7'h64 == i ? a_100 : _GEN_99;
  assign _GEN_101 = 7'h65 == i ? a_101 : _GEN_100;
  assign _GEN_102 = 7'h66 == i ? a_102 : _GEN_101;
  assign _GEN_103 = 7'h67 == i ? a_103 : _GEN_102;
  assign _GEN_104 = 7'h68 == i ? a_104 : _GEN_103;
  assign _GEN_105 = 7'h69 == i ? a_105 : _GEN_104;
  assign _GEN_106 = 7'h6a == i ? a_106 : _GEN_105;
  assign _GEN_107 = 7'h6b == i ? a_107 : _GEN_106;
  assign _GEN_108 = 7'h6c == i ? a_108 : _GEN_107;
  assign _GEN_109 = 7'h6d == i ? a_109 : _GEN_108;
  assign _GEN_110 = 7'h6e == i ? a_110 : _GEN_109;
  assign _GEN_111 = 7'h6f == i ? a_111 : _GEN_110;
  assign _GEN_112 = 7'h70 == i ? a_112 : _GEN_111;
  assign _GEN_113 = 7'h71 == i ? a_113 : _GEN_112;
  assign _GEN_114 = 7'h72 == i ? a_114 : _GEN_113;
  assign _GEN_115 = 7'h73 == i ? a_115 : _GEN_114;
  assign _GEN_116 = 7'h74 == i ? a_116 : _GEN_115;
  assign _GEN_117 = 7'h75 == i ? a_117 : _GEN_116;
  assign _GEN_118 = 7'h76 == i ? a_118 : _GEN_117;
  assign _GEN_119 = 7'h77 == i ? a_119 : _GEN_118;
  assign _GEN_121 = 7'h1 == i ? b_1 : b_0;
  assign _GEN_122 = 7'h2 == i ? b_2 : _GEN_121;
  assign _GEN_123 = 7'h3 == i ? b_3 : _GEN_122;
  assign _GEN_124 = 7'h4 == i ? b_4 : _GEN_123;
  assign _GEN_125 = 7'h5 == i ? b_5 : _GEN_124;
  assign _GEN_126 = 7'h6 == i ? b_6 : _GEN_125;
  assign _GEN_127 = 7'h7 == i ? b_7 : _GEN_126;
  assign _GEN_128 = 7'h8 == i ? b_8 : _GEN_127;
  assign _GEN_129 = 7'h9 == i ? b_9 : _GEN_128;
  assign _GEN_130 = 7'ha == i ? b_10 : _GEN_129;
  assign _GEN_131 = 7'hb == i ? b_11 : _GEN_130;
  assign _GEN_132 = 7'hc == i ? b_12 : _GEN_131;
  assign _GEN_133 = 7'hd == i ? b_13 : _GEN_132;
  assign _GEN_134 = 7'he == i ? b_14 : _GEN_133;
  assign _GEN_135 = 7'hf == i ? b_15 : _GEN_134;
  assign _GEN_136 = 7'h10 == i ? b_16 : _GEN_135;
  assign _GEN_137 = 7'h11 == i ? b_17 : _GEN_136;
  assign _GEN_138 = 7'h12 == i ? b_18 : _GEN_137;
  assign _GEN_139 = 7'h13 == i ? b_19 : _GEN_138;
  assign _GEN_140 = 7'h14 == i ? b_20 : _GEN_139;
  assign _GEN_141 = 7'h15 == i ? b_21 : _GEN_140;
  assign _GEN_142 = 7'h16 == i ? b_22 : _GEN_141;
  assign _GEN_143 = 7'h17 == i ? b_23 : _GEN_142;
  assign _GEN_144 = 7'h18 == i ? b_24 : _GEN_143;
  assign _GEN_145 = 7'h19 == i ? b_25 : _GEN_144;
  assign _GEN_146 = 7'h1a == i ? b_26 : _GEN_145;
  assign _GEN_147 = 7'h1b == i ? b_27 : _GEN_146;
  assign _GEN_148 = 7'h1c == i ? b_28 : _GEN_147;
  assign _GEN_149 = 7'h1d == i ? b_29 : _GEN_148;
  assign _GEN_150 = 7'h1e == i ? b_30 : _GEN_149;
  assign _GEN_151 = 7'h1f == i ? b_31 : _GEN_150;
  assign _GEN_152 = 7'h20 == i ? b_32 : _GEN_151;
  assign _GEN_153 = 7'h21 == i ? b_33 : _GEN_152;
  assign _GEN_154 = 7'h22 == i ? b_34 : _GEN_153;
  assign _GEN_155 = 7'h23 == i ? b_35 : _GEN_154;
  assign _GEN_156 = 7'h24 == i ? b_36 : _GEN_155;
  assign _GEN_157 = 7'h25 == i ? b_37 : _GEN_156;
  assign _GEN_158 = 7'h26 == i ? b_38 : _GEN_157;
  assign _GEN_159 = 7'h27 == i ? b_39 : _GEN_158;
  assign _GEN_160 = 7'h28 == i ? b_40 : _GEN_159;
  assign _GEN_161 = 7'h29 == i ? b_41 : _GEN_160;
  assign _GEN_162 = 7'h2a == i ? b_42 : _GEN_161;
  assign _GEN_163 = 7'h2b == i ? b_43 : _GEN_162;
  assign _GEN_164 = 7'h2c == i ? b_44 : _GEN_163;
  assign _GEN_165 = 7'h2d == i ? b_45 : _GEN_164;
  assign _GEN_166 = 7'h2e == i ? b_46 : _GEN_165;
  assign _GEN_167 = 7'h2f == i ? b_47 : _GEN_166;
  assign _GEN_168 = 7'h30 == i ? b_48 : _GEN_167;
  assign _GEN_169 = 7'h31 == i ? b_49 : _GEN_168;
  assign _GEN_170 = 7'h32 == i ? b_50 : _GEN_169;
  assign _GEN_171 = 7'h33 == i ? b_51 : _GEN_170;
  assign _GEN_172 = 7'h34 == i ? b_52 : _GEN_171;
  assign _GEN_173 = 7'h35 == i ? b_53 : _GEN_172;
  assign _GEN_174 = 7'h36 == i ? b_54 : _GEN_173;
  assign _GEN_175 = 7'h37 == i ? b_55 : _GEN_174;
  assign _GEN_176 = 7'h38 == i ? b_56 : _GEN_175;
  assign _GEN_177 = 7'h39 == i ? b_57 : _GEN_176;
  assign _GEN_178 = 7'h3a == i ? b_58 : _GEN_177;
  assign _GEN_179 = 7'h3b == i ? b_59 : _GEN_178;
  assign _GEN_180 = 7'h3c == i ? b_60 : _GEN_179;
  assign _GEN_181 = 7'h3d == i ? b_61 : _GEN_180;
  assign _GEN_182 = 7'h3e == i ? b_62 : _GEN_181;
  assign _GEN_183 = 7'h3f == i ? b_63 : _GEN_182;
  assign _GEN_184 = 7'h40 == i ? b_64 : _GEN_183;
  assign _GEN_185 = 7'h41 == i ? b_65 : _GEN_184;
  assign _GEN_186 = 7'h42 == i ? b_66 : _GEN_185;
  assign _GEN_187 = 7'h43 == i ? b_67 : _GEN_186;
  assign _GEN_188 = 7'h44 == i ? b_68 : _GEN_187;
  assign _GEN_189 = 7'h45 == i ? b_69 : _GEN_188;
  assign _GEN_190 = 7'h46 == i ? b_70 : _GEN_189;
  assign _GEN_191 = 7'h47 == i ? b_71 : _GEN_190;
  assign _GEN_192 = 7'h48 == i ? b_72 : _GEN_191;
  assign _GEN_193 = 7'h49 == i ? b_73 : _GEN_192;
  assign _GEN_194 = 7'h4a == i ? b_74 : _GEN_193;
  assign _GEN_195 = 7'h4b == i ? b_75 : _GEN_194;
  assign _GEN_196 = 7'h4c == i ? b_76 : _GEN_195;
  assign _GEN_197 = 7'h4d == i ? b_77 : _GEN_196;
  assign _GEN_198 = 7'h4e == i ? b_78 : _GEN_197;
  assign _GEN_199 = 7'h4f == i ? b_79 : _GEN_198;
  assign _GEN_200 = 7'h50 == i ? b_80 : _GEN_199;
  assign _GEN_201 = 7'h51 == i ? b_81 : _GEN_200;
  assign _GEN_202 = 7'h52 == i ? b_82 : _GEN_201;
  assign _GEN_203 = 7'h53 == i ? b_83 : _GEN_202;
  assign _GEN_204 = 7'h54 == i ? b_84 : _GEN_203;
  assign _GEN_205 = 7'h55 == i ? b_85 : _GEN_204;
  assign _GEN_206 = 7'h56 == i ? b_86 : _GEN_205;
  assign _GEN_207 = 7'h57 == i ? b_87 : _GEN_206;
  assign _GEN_208 = 7'h58 == i ? b_88 : _GEN_207;
  assign _GEN_209 = 7'h59 == i ? b_89 : _GEN_208;
  assign _GEN_210 = 7'h5a == i ? b_90 : _GEN_209;
  assign _GEN_211 = 7'h5b == i ? b_91 : _GEN_210;
  assign _GEN_212 = 7'h5c == i ? b_92 : _GEN_211;
  assign _GEN_213 = 7'h5d == i ? b_93 : _GEN_212;
  assign _GEN_214 = 7'h5e == i ? b_94 : _GEN_213;
  assign _GEN_215 = 7'h5f == i ? b_95 : _GEN_214;
  assign _GEN_216 = 7'h60 == i ? b_96 : _GEN_215;
  assign _GEN_217 = 7'h61 == i ? b_97 : _GEN_216;
  assign _GEN_218 = 7'h62 == i ? b_98 : _GEN_217;
  assign _GEN_219 = 7'h63 == i ? b_99 : _GEN_218;
  assign _GEN_220 = 7'h64 == i ? b_100 : _GEN_219;
  assign _GEN_221 = 7'h65 == i ? b_101 : _GEN_220;
  assign _GEN_222 = 7'h66 == i ? b_102 : _GEN_221;
  assign _GEN_223 = 7'h67 == i ? b_103 : _GEN_222;
  assign _GEN_224 = 7'h68 == i ? b_104 : _GEN_223;
  assign _GEN_225 = 7'h69 == i ? b_105 : _GEN_224;
  assign _GEN_226 = 7'h6a == i ? b_106 : _GEN_225;
  assign _GEN_227 = 7'h6b == i ? b_107 : _GEN_226;
  assign _GEN_228 = 7'h6c == i ? b_108 : _GEN_227;
  assign _GEN_229 = 7'h6d == i ? b_109 : _GEN_228;
  assign _GEN_230 = 7'h6e == i ? b_110 : _GEN_229;
  assign _GEN_231 = 7'h6f == i ? b_111 : _GEN_230;
  assign _GEN_232 = 7'h70 == i ? b_112 : _GEN_231;
  assign _GEN_233 = 7'h71 == i ? b_113 : _GEN_232;
  assign _GEN_234 = 7'h72 == i ? b_114 : _GEN_233;
  assign _GEN_235 = 7'h73 == i ? b_115 : _GEN_234;
  assign _GEN_236 = 7'h74 == i ? b_116 : _GEN_235;
  assign _GEN_237 = 7'h75 == i ? b_117 : _GEN_236;
  assign _GEN_238 = 7'h76 == i ? b_118 : _GEN_237;
  assign _GEN_239 = 7'h77 == i ? b_119 : _GEN_238;
  assign _T_240 = _GEN_119 * _GEN_239;
  assign _T_241 = sum + _T_240;
  assign _T_242 = i + 7'h1;
  assign _GEN_240 = _T_244 ? _T_242 : 8'h0;
  assign _GEN_241 = _T_244 ? _T_241 : 33'h0;
  assign _GEN_242 = _T_243 ? 8'h0 : _GEN_240;
  assign _GEN_244 = _T_243 ? sum : 32'h0;
  assign _GEN_245 = _T_243 ? 33'h0 : _GEN_241;
  assign _GEN_246 = io_rdy ? _T_241 : _GEN_245;
  assign _GEN_247 = io_rdy ? _T_242 : _GEN_242;
  assign io_q = io_rdy ? 32'h0 : _GEN_244;
  assign io_v = io_rdy ? 1'h0 : _T_243;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sum = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  i = _RAND_1[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      sum <= 32'h0;
    end else begin
      sum <= _GEN_246[31:0];
    end
    if (reset) begin
      i <= 7'h0;
    end else begin
      i <= _GEN_247[6:0];
    end
  end
endmodule
module Node_103(
  input           clock,
  input           reset,
  input  [1919:0] io_d_in,
  input  [1919:0] io_w,
  input           io_rdy,
  input  [15:0]   io_bias,
  output [15:0]   io_d_out,
  output          io_v
);
  wire  muladdc_clock;
  wire  muladdc_reset;
  wire [1919:0] muladdc_io_a;
  wire [1919:0] muladdc_io_b;
  wire  muladdc_io_rdy;
  wire [31:0] muladdc_io_q;
  wire  muladdc_io_v;
  wire [31:0] act_io_q;
  wire [15:0] act_io_bias;
  wire  act_io_v_in;
  wire [15:0] act_io_d;
  wire  act_io_v_out;
  Mac_103 muladdc (
    .clock(muladdc_clock),
    .reset(muladdc_reset),
    .io_a(muladdc_io_a),
    .io_b(muladdc_io_b),
    .io_rdy(muladdc_io_rdy),
    .io_q(muladdc_io_q),
    .io_v(muladdc_io_v)
  );
  ReLU act (
    .io_q(act_io_q),
    .io_bias(act_io_bias),
    .io_v_in(act_io_v_in),
    .io_d(act_io_d),
    .io_v_out(act_io_v_out)
  );
  assign io_d_out = act_io_d;
  assign io_v = act_io_v_out;
  assign muladdc_clock = clock;
  assign muladdc_reset = reset;
  assign muladdc_io_a = io_d_in;
  assign muladdc_io_b = io_w;
  assign muladdc_io_rdy = io_rdy;
  assign act_io_q = muladdc_io_q;
  assign act_io_bias = io_bias;
  assign act_io_v_in = muladdc_io_v;
endmodule
module FC2(
  input           clock,
  input           reset,
  input  [15:0]   io_d_in,
  input  [1919:0] io_w_in,
  input  [15:0]   io_bias,
  input           io_rdy,
  input           io_done,
  output [15:0]   io_d_out,
  output          io_v,
  output          io_fc1_done
);
  wire  in_channel_clock;
  wire  in_channel_reset;
  wire [15:0] in_channel_io_d_in;
  wire  in_channel_io_en;
  wire [1919:0] in_channel_io_d_out;
  wire  conv_node2_clock;
  wire  conv_node2_reset;
  wire [1919:0] conv_node2_io_d_in;
  wire [1919:0] conv_node2_io_w;
  wire  conv_node2_io_rdy;
  wire [15:0] conv_node2_io_bias;
  wire [15:0] conv_node2_io_d_out;
  wire  conv_node2_io_v;
  reg  rdy;
  reg [31:0] _RAND_0;
  reg [1919:0] store;
  reg [1919:0] _RAND_1;
  reg  first_rdy;
  reg [31:0] _RAND_2;
  reg [15:0] in_counter;
  reg [31:0] _RAND_3;
  wire  _T;
  wire [16:0] _T_1;
  wire [16:0] _GEN_0;
  wire [16:0] _GEN_1;
  reg  is_done;
  reg [31:0] _RAND_4;
  wire  _GEN_4;
  wire  _T_2;
  ShiftRegister_22 in_channel (
    .clock(in_channel_clock),
    .reset(in_channel_reset),
    .io_d_in(in_channel_io_d_in),
    .io_en(in_channel_io_en),
    .io_d_out(in_channel_io_d_out)
  );
  Node_103 conv_node2 (
    .clock(conv_node2_clock),
    .reset(conv_node2_reset),
    .io_d_in(conv_node2_io_d_in),
    .io_w(conv_node2_io_w),
    .io_rdy(conv_node2_io_rdy),
    .io_bias(conv_node2_io_bias),
    .io_d_out(conv_node2_io_d_out),
    .io_v(conv_node2_io_v)
  );
  assign _T = in_counter == 16'h78;
  assign _T_1 = in_counter + 16'h1;
  assign _GEN_0 = io_rdy ? _T_1 : {{1'd0}, in_counter};
  assign _GEN_1 = _T ? 17'h0 : _GEN_0;
  assign _GEN_4 = io_done | is_done;
  assign _T_2 = first_rdy | conv_node2_io_v;
  assign io_d_out = conv_node2_io_d_out;
  assign io_v = conv_node2_io_v;
  assign io_fc1_done = in_counter == 16'h78;
  assign in_channel_clock = clock;
  assign in_channel_reset = reset;
  assign in_channel_io_d_in = io_d_in;
  assign in_channel_io_en = io_rdy;
  assign conv_node2_clock = clock;
  assign conv_node2_reset = reset;
  assign conv_node2_io_d_in = store;
  assign conv_node2_io_w = io_w_in;
  assign conv_node2_io_rdy = rdy;
  assign conv_node2_io_bias = io_bias;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rdy = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {60{`RANDOM}};
  store = _RAND_1[1919:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  first_rdy = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_counter = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  is_done = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      rdy <= 1'h0;
    end else if (is_done) begin
      rdy <= 1'h0;
    end else begin
      rdy <= _T_2;
    end
    if (reset) begin
      store <= 1920'h0;
    end else if (_T) begin
      store <= in_channel_io_d_out;
    end
    if (reset) begin
      first_rdy <= 1'h0;
    end else begin
      first_rdy <= _T;
    end
    if (reset) begin
      in_counter <= 16'h0;
    end else begin
      in_counter <= _GEN_1[15:0];
    end
    if (reset) begin
      is_done <= 1'h0;
    end else begin
      is_done <= _GEN_4;
    end
  end
endmodule
module ShiftRegister_23(
  input           clock,
  input           reset,
  input  [15:0]   io_d_in,
  input           io_en,
  output [1343:0] io_d_out
);
  reg [15:0] _T;
  reg [31:0] _RAND_0;
  reg [15:0] _T_1;
  reg [31:0] _RAND_1;
  reg [15:0] _T_2;
  reg [31:0] _RAND_2;
  reg [15:0] _T_3;
  reg [31:0] _RAND_3;
  reg [15:0] _T_4;
  reg [31:0] _RAND_4;
  reg [15:0] _T_5;
  reg [31:0] _RAND_5;
  reg [15:0] _T_6;
  reg [31:0] _RAND_6;
  reg [15:0] _T_7;
  reg [31:0] _RAND_7;
  reg [15:0] _T_8;
  reg [31:0] _RAND_8;
  reg [15:0] _T_9;
  reg [31:0] _RAND_9;
  reg [15:0] _T_10;
  reg [31:0] _RAND_10;
  reg [15:0] _T_11;
  reg [31:0] _RAND_11;
  reg [15:0] _T_12;
  reg [31:0] _RAND_12;
  reg [15:0] _T_13;
  reg [31:0] _RAND_13;
  reg [15:0] _T_14;
  reg [31:0] _RAND_14;
  reg [15:0] _T_15;
  reg [31:0] _RAND_15;
  reg [15:0] _T_16;
  reg [31:0] _RAND_16;
  reg [15:0] _T_17;
  reg [31:0] _RAND_17;
  reg [15:0] _T_18;
  reg [31:0] _RAND_18;
  reg [15:0] _T_19;
  reg [31:0] _RAND_19;
  reg [15:0] _T_20;
  reg [31:0] _RAND_20;
  reg [15:0] _T_21;
  reg [31:0] _RAND_21;
  reg [15:0] _T_22;
  reg [31:0] _RAND_22;
  reg [15:0] _T_23;
  reg [31:0] _RAND_23;
  reg [15:0] _T_24;
  reg [31:0] _RAND_24;
  reg [15:0] _T_25;
  reg [31:0] _RAND_25;
  reg [15:0] _T_26;
  reg [31:0] _RAND_26;
  reg [15:0] _T_27;
  reg [31:0] _RAND_27;
  reg [15:0] _T_28;
  reg [31:0] _RAND_28;
  reg [15:0] _T_29;
  reg [31:0] _RAND_29;
  reg [15:0] _T_30;
  reg [31:0] _RAND_30;
  reg [15:0] _T_31;
  reg [31:0] _RAND_31;
  reg [15:0] _T_32;
  reg [31:0] _RAND_32;
  reg [15:0] _T_33;
  reg [31:0] _RAND_33;
  reg [15:0] _T_34;
  reg [31:0] _RAND_34;
  reg [15:0] _T_35;
  reg [31:0] _RAND_35;
  reg [15:0] _T_36;
  reg [31:0] _RAND_36;
  reg [15:0] _T_37;
  reg [31:0] _RAND_37;
  reg [15:0] _T_38;
  reg [31:0] _RAND_38;
  reg [15:0] _T_39;
  reg [31:0] _RAND_39;
  reg [15:0] _T_40;
  reg [31:0] _RAND_40;
  reg [15:0] _T_41;
  reg [31:0] _RAND_41;
  reg [15:0] _T_42;
  reg [31:0] _RAND_42;
  reg [15:0] _T_43;
  reg [31:0] _RAND_43;
  reg [15:0] _T_44;
  reg [31:0] _RAND_44;
  reg [15:0] _T_45;
  reg [31:0] _RAND_45;
  reg [15:0] _T_46;
  reg [31:0] _RAND_46;
  reg [15:0] _T_47;
  reg [31:0] _RAND_47;
  reg [15:0] _T_48;
  reg [31:0] _RAND_48;
  reg [15:0] _T_49;
  reg [31:0] _RAND_49;
  reg [15:0] _T_50;
  reg [31:0] _RAND_50;
  reg [15:0] _T_51;
  reg [31:0] _RAND_51;
  reg [15:0] _T_52;
  reg [31:0] _RAND_52;
  reg [15:0] _T_53;
  reg [31:0] _RAND_53;
  reg [15:0] _T_54;
  reg [31:0] _RAND_54;
  reg [15:0] _T_55;
  reg [31:0] _RAND_55;
  reg [15:0] _T_56;
  reg [31:0] _RAND_56;
  reg [15:0] _T_57;
  reg [31:0] _RAND_57;
  reg [15:0] _T_58;
  reg [31:0] _RAND_58;
  reg [15:0] _T_59;
  reg [31:0] _RAND_59;
  reg [15:0] _T_60;
  reg [31:0] _RAND_60;
  reg [15:0] _T_61;
  reg [31:0] _RAND_61;
  reg [15:0] _T_62;
  reg [31:0] _RAND_62;
  reg [15:0] _T_63;
  reg [31:0] _RAND_63;
  reg [15:0] _T_64;
  reg [31:0] _RAND_64;
  reg [15:0] _T_65;
  reg [31:0] _RAND_65;
  reg [15:0] _T_66;
  reg [31:0] _RAND_66;
  reg [15:0] _T_67;
  reg [31:0] _RAND_67;
  reg [15:0] _T_68;
  reg [31:0] _RAND_68;
  reg [15:0] _T_69;
  reg [31:0] _RAND_69;
  reg [15:0] _T_70;
  reg [31:0] _RAND_70;
  reg [15:0] _T_71;
  reg [31:0] _RAND_71;
  reg [15:0] _T_72;
  reg [31:0] _RAND_72;
  reg [15:0] _T_73;
  reg [31:0] _RAND_73;
  reg [15:0] _T_74;
  reg [31:0] _RAND_74;
  reg [15:0] _T_75;
  reg [31:0] _RAND_75;
  reg [15:0] _T_76;
  reg [31:0] _RAND_76;
  reg [15:0] _T_77;
  reg [31:0] _RAND_77;
  reg [15:0] _T_78;
  reg [31:0] _RAND_78;
  reg [15:0] _T_79;
  reg [31:0] _RAND_79;
  reg [15:0] _T_80;
  reg [31:0] _RAND_80;
  reg [15:0] _T_81;
  reg [31:0] _RAND_81;
  reg [15:0] _T_82;
  reg [31:0] _RAND_82;
  reg [15:0] _T_83;
  reg [31:0] _RAND_83;
  wire [159:0] _T_92;
  wire [95:0] _T_101;
  wire [159:0] _T_112;
  wire [95:0] _T_121;
  wire [335:0] _T_123;
  wire [671:0] _T_124;
  wire [159:0] _T_133;
  wire [95:0] _T_142;
  wire [159:0] _T_153;
  wire [95:0] _T_162;
  wire [335:0] _T_164;
  wire [671:0] _T_165;
  assign _T_92 = {_T,_T_1,_T_2,_T_3,_T_4,_T_5,_T_6,_T_7,_T_8,_T_9};
  assign _T_101 = {_T_15,_T_16,_T_17,_T_18,_T_19,_T_20};
  assign _T_112 = {_T_21,_T_22,_T_23,_T_24,_T_25,_T_26,_T_27,_T_28,_T_29,_T_30};
  assign _T_121 = {_T_36,_T_37,_T_38,_T_39,_T_40,_T_41};
  assign _T_123 = {_T_112,_T_31,_T_32,_T_33,_T_34,_T_35,_T_121};
  assign _T_124 = {_T_92,_T_10,_T_11,_T_12,_T_13,_T_14,_T_101,_T_123};
  assign _T_133 = {_T_42,_T_43,_T_44,_T_45,_T_46,_T_47,_T_48,_T_49,_T_50,_T_51};
  assign _T_142 = {_T_57,_T_58,_T_59,_T_60,_T_61,_T_62};
  assign _T_153 = {_T_63,_T_64,_T_65,_T_66,_T_67,_T_68,_T_69,_T_70,_T_71,_T_72};
  assign _T_162 = {_T_78,_T_79,_T_80,_T_81,_T_82,_T_83};
  assign _T_164 = {_T_153,_T_73,_T_74,_T_75,_T_76,_T_77,_T_162};
  assign _T_165 = {_T_133,_T_52,_T_53,_T_54,_T_55,_T_56,_T_142,_T_164};
  assign io_d_out = {_T_124,_T_165};
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_6 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_7 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_8 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_9 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_10 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_11 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_12 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_13 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_14 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_15 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_16 = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_17 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_18 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_19 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_20 = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_21 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_22 = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_23 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_24 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_25 = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_26 = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_27 = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_28 = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_29 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_30 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_31 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_32 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_33 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_34 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_35 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_36 = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_37 = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_38 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_39 = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_40 = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_41 = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_42 = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_43 = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_44 = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_45 = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_46 = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_47 = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_48 = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_49 = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_50 = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_51 = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_52 = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_53 = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_54 = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_55 = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_56 = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_57 = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_58 = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_59 = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_60 = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_61 = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_62 = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_63 = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_64 = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_65 = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_66 = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_67 = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_68 = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_69 = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_70 = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_71 = _RAND_71[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_72 = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_73 = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_74 = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_75 = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_76 = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_77 = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_78 = _RAND_78[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_79 = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_80 = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_81 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_82 = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_83 = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T <= 16'h0;
    end else if (io_en) begin
      _T <= io_d_in;
    end
    if (reset) begin
      _T_1 <= 16'h0;
    end else if (io_en) begin
      _T_1 <= _T;
    end
    if (reset) begin
      _T_2 <= 16'h0;
    end else if (io_en) begin
      _T_2 <= _T_1;
    end
    if (reset) begin
      _T_3 <= 16'h0;
    end else if (io_en) begin
      _T_3 <= _T_2;
    end
    if (reset) begin
      _T_4 <= 16'h0;
    end else if (io_en) begin
      _T_4 <= _T_3;
    end
    if (reset) begin
      _T_5 <= 16'h0;
    end else if (io_en) begin
      _T_5 <= _T_4;
    end
    if (reset) begin
      _T_6 <= 16'h0;
    end else if (io_en) begin
      _T_6 <= _T_5;
    end
    if (reset) begin
      _T_7 <= 16'h0;
    end else if (io_en) begin
      _T_7 <= _T_6;
    end
    if (reset) begin
      _T_8 <= 16'h0;
    end else if (io_en) begin
      _T_8 <= _T_7;
    end
    if (reset) begin
      _T_9 <= 16'h0;
    end else if (io_en) begin
      _T_9 <= _T_8;
    end
    if (reset) begin
      _T_10 <= 16'h0;
    end else if (io_en) begin
      _T_10 <= _T_9;
    end
    if (reset) begin
      _T_11 <= 16'h0;
    end else if (io_en) begin
      _T_11 <= _T_10;
    end
    if (reset) begin
      _T_12 <= 16'h0;
    end else if (io_en) begin
      _T_12 <= _T_11;
    end
    if (reset) begin
      _T_13 <= 16'h0;
    end else if (io_en) begin
      _T_13 <= _T_12;
    end
    if (reset) begin
      _T_14 <= 16'h0;
    end else if (io_en) begin
      _T_14 <= _T_13;
    end
    if (reset) begin
      _T_15 <= 16'h0;
    end else if (io_en) begin
      _T_15 <= _T_14;
    end
    if (reset) begin
      _T_16 <= 16'h0;
    end else if (io_en) begin
      _T_16 <= _T_15;
    end
    if (reset) begin
      _T_17 <= 16'h0;
    end else if (io_en) begin
      _T_17 <= _T_16;
    end
    if (reset) begin
      _T_18 <= 16'h0;
    end else if (io_en) begin
      _T_18 <= _T_17;
    end
    if (reset) begin
      _T_19 <= 16'h0;
    end else if (io_en) begin
      _T_19 <= _T_18;
    end
    if (reset) begin
      _T_20 <= 16'h0;
    end else if (io_en) begin
      _T_20 <= _T_19;
    end
    if (reset) begin
      _T_21 <= 16'h0;
    end else if (io_en) begin
      _T_21 <= _T_20;
    end
    if (reset) begin
      _T_22 <= 16'h0;
    end else if (io_en) begin
      _T_22 <= _T_21;
    end
    if (reset) begin
      _T_23 <= 16'h0;
    end else if (io_en) begin
      _T_23 <= _T_22;
    end
    if (reset) begin
      _T_24 <= 16'h0;
    end else if (io_en) begin
      _T_24 <= _T_23;
    end
    if (reset) begin
      _T_25 <= 16'h0;
    end else if (io_en) begin
      _T_25 <= _T_24;
    end
    if (reset) begin
      _T_26 <= 16'h0;
    end else if (io_en) begin
      _T_26 <= _T_25;
    end
    if (reset) begin
      _T_27 <= 16'h0;
    end else if (io_en) begin
      _T_27 <= _T_26;
    end
    if (reset) begin
      _T_28 <= 16'h0;
    end else if (io_en) begin
      _T_28 <= _T_27;
    end
    if (reset) begin
      _T_29 <= 16'h0;
    end else if (io_en) begin
      _T_29 <= _T_28;
    end
    if (reset) begin
      _T_30 <= 16'h0;
    end else if (io_en) begin
      _T_30 <= _T_29;
    end
    if (reset) begin
      _T_31 <= 16'h0;
    end else if (io_en) begin
      _T_31 <= _T_30;
    end
    if (reset) begin
      _T_32 <= 16'h0;
    end else if (io_en) begin
      _T_32 <= _T_31;
    end
    if (reset) begin
      _T_33 <= 16'h0;
    end else if (io_en) begin
      _T_33 <= _T_32;
    end
    if (reset) begin
      _T_34 <= 16'h0;
    end else if (io_en) begin
      _T_34 <= _T_33;
    end
    if (reset) begin
      _T_35 <= 16'h0;
    end else if (io_en) begin
      _T_35 <= _T_34;
    end
    if (reset) begin
      _T_36 <= 16'h0;
    end else if (io_en) begin
      _T_36 <= _T_35;
    end
    if (reset) begin
      _T_37 <= 16'h0;
    end else if (io_en) begin
      _T_37 <= _T_36;
    end
    if (reset) begin
      _T_38 <= 16'h0;
    end else if (io_en) begin
      _T_38 <= _T_37;
    end
    if (reset) begin
      _T_39 <= 16'h0;
    end else if (io_en) begin
      _T_39 <= _T_38;
    end
    if (reset) begin
      _T_40 <= 16'h0;
    end else if (io_en) begin
      _T_40 <= _T_39;
    end
    if (reset) begin
      _T_41 <= 16'h0;
    end else if (io_en) begin
      _T_41 <= _T_40;
    end
    if (reset) begin
      _T_42 <= 16'h0;
    end else if (io_en) begin
      _T_42 <= _T_41;
    end
    if (reset) begin
      _T_43 <= 16'h0;
    end else if (io_en) begin
      _T_43 <= _T_42;
    end
    if (reset) begin
      _T_44 <= 16'h0;
    end else if (io_en) begin
      _T_44 <= _T_43;
    end
    if (reset) begin
      _T_45 <= 16'h0;
    end else if (io_en) begin
      _T_45 <= _T_44;
    end
    if (reset) begin
      _T_46 <= 16'h0;
    end else if (io_en) begin
      _T_46 <= _T_45;
    end
    if (reset) begin
      _T_47 <= 16'h0;
    end else if (io_en) begin
      _T_47 <= _T_46;
    end
    if (reset) begin
      _T_48 <= 16'h0;
    end else if (io_en) begin
      _T_48 <= _T_47;
    end
    if (reset) begin
      _T_49 <= 16'h0;
    end else if (io_en) begin
      _T_49 <= _T_48;
    end
    if (reset) begin
      _T_50 <= 16'h0;
    end else if (io_en) begin
      _T_50 <= _T_49;
    end
    if (reset) begin
      _T_51 <= 16'h0;
    end else if (io_en) begin
      _T_51 <= _T_50;
    end
    if (reset) begin
      _T_52 <= 16'h0;
    end else if (io_en) begin
      _T_52 <= _T_51;
    end
    if (reset) begin
      _T_53 <= 16'h0;
    end else if (io_en) begin
      _T_53 <= _T_52;
    end
    if (reset) begin
      _T_54 <= 16'h0;
    end else if (io_en) begin
      _T_54 <= _T_53;
    end
    if (reset) begin
      _T_55 <= 16'h0;
    end else if (io_en) begin
      _T_55 <= _T_54;
    end
    if (reset) begin
      _T_56 <= 16'h0;
    end else if (io_en) begin
      _T_56 <= _T_55;
    end
    if (reset) begin
      _T_57 <= 16'h0;
    end else if (io_en) begin
      _T_57 <= _T_56;
    end
    if (reset) begin
      _T_58 <= 16'h0;
    end else if (io_en) begin
      _T_58 <= _T_57;
    end
    if (reset) begin
      _T_59 <= 16'h0;
    end else if (io_en) begin
      _T_59 <= _T_58;
    end
    if (reset) begin
      _T_60 <= 16'h0;
    end else if (io_en) begin
      _T_60 <= _T_59;
    end
    if (reset) begin
      _T_61 <= 16'h0;
    end else if (io_en) begin
      _T_61 <= _T_60;
    end
    if (reset) begin
      _T_62 <= 16'h0;
    end else if (io_en) begin
      _T_62 <= _T_61;
    end
    if (reset) begin
      _T_63 <= 16'h0;
    end else if (io_en) begin
      _T_63 <= _T_62;
    end
    if (reset) begin
      _T_64 <= 16'h0;
    end else if (io_en) begin
      _T_64 <= _T_63;
    end
    if (reset) begin
      _T_65 <= 16'h0;
    end else if (io_en) begin
      _T_65 <= _T_64;
    end
    if (reset) begin
      _T_66 <= 16'h0;
    end else if (io_en) begin
      _T_66 <= _T_65;
    end
    if (reset) begin
      _T_67 <= 16'h0;
    end else if (io_en) begin
      _T_67 <= _T_66;
    end
    if (reset) begin
      _T_68 <= 16'h0;
    end else if (io_en) begin
      _T_68 <= _T_67;
    end
    if (reset) begin
      _T_69 <= 16'h0;
    end else if (io_en) begin
      _T_69 <= _T_68;
    end
    if (reset) begin
      _T_70 <= 16'h0;
    end else if (io_en) begin
      _T_70 <= _T_69;
    end
    if (reset) begin
      _T_71 <= 16'h0;
    end else if (io_en) begin
      _T_71 <= _T_70;
    end
    if (reset) begin
      _T_72 <= 16'h0;
    end else if (io_en) begin
      _T_72 <= _T_71;
    end
    if (reset) begin
      _T_73 <= 16'h0;
    end else if (io_en) begin
      _T_73 <= _T_72;
    end
    if (reset) begin
      _T_74 <= 16'h0;
    end else if (io_en) begin
      _T_74 <= _T_73;
    end
    if (reset) begin
      _T_75 <= 16'h0;
    end else if (io_en) begin
      _T_75 <= _T_74;
    end
    if (reset) begin
      _T_76 <= 16'h0;
    end else if (io_en) begin
      _T_76 <= _T_75;
    end
    if (reset) begin
      _T_77 <= 16'h0;
    end else if (io_en) begin
      _T_77 <= _T_76;
    end
    if (reset) begin
      _T_78 <= 16'h0;
    end else if (io_en) begin
      _T_78 <= _T_77;
    end
    if (reset) begin
      _T_79 <= 16'h0;
    end else if (io_en) begin
      _T_79 <= _T_78;
    end
    if (reset) begin
      _T_80 <= 16'h0;
    end else if (io_en) begin
      _T_80 <= _T_79;
    end
    if (reset) begin
      _T_81 <= 16'h0;
    end else if (io_en) begin
      _T_81 <= _T_80;
    end
    if (reset) begin
      _T_82 <= 16'h0;
    end else if (io_en) begin
      _T_82 <= _T_81;
    end
    if (reset) begin
      _T_83 <= 16'h0;
    end else if (io_en) begin
      _T_83 <= _T_82;
    end
  end
endmodule
module Mac_104(
  input           clock,
  input           reset,
  input  [1343:0] io_a,
  input  [1343:0] io_b,
  input           io_rdy,
  output [31:0]   io_q,
  output          io_v
);
  wire [15:0] a_0;
  wire [15:0] b_0;
  wire [15:0] a_1;
  wire [15:0] b_1;
  wire [15:0] a_2;
  wire [15:0] b_2;
  wire [15:0] a_3;
  wire [15:0] b_3;
  wire [15:0] a_4;
  wire [15:0] b_4;
  wire [15:0] a_5;
  wire [15:0] b_5;
  wire [15:0] a_6;
  wire [15:0] b_6;
  wire [15:0] a_7;
  wire [15:0] b_7;
  wire [15:0] a_8;
  wire [15:0] b_8;
  wire [15:0] a_9;
  wire [15:0] b_9;
  wire [15:0] a_10;
  wire [15:0] b_10;
  wire [15:0] a_11;
  wire [15:0] b_11;
  wire [15:0] a_12;
  wire [15:0] b_12;
  wire [15:0] a_13;
  wire [15:0] b_13;
  wire [15:0] a_14;
  wire [15:0] b_14;
  wire [15:0] a_15;
  wire [15:0] b_15;
  wire [15:0] a_16;
  wire [15:0] b_16;
  wire [15:0] a_17;
  wire [15:0] b_17;
  wire [15:0] a_18;
  wire [15:0] b_18;
  wire [15:0] a_19;
  wire [15:0] b_19;
  wire [15:0] a_20;
  wire [15:0] b_20;
  wire [15:0] a_21;
  wire [15:0] b_21;
  wire [15:0] a_22;
  wire [15:0] b_22;
  wire [15:0] a_23;
  wire [15:0] b_23;
  wire [15:0] a_24;
  wire [15:0] b_24;
  wire [15:0] a_25;
  wire [15:0] b_25;
  wire [15:0] a_26;
  wire [15:0] b_26;
  wire [15:0] a_27;
  wire [15:0] b_27;
  wire [15:0] a_28;
  wire [15:0] b_28;
  wire [15:0] a_29;
  wire [15:0] b_29;
  wire [15:0] a_30;
  wire [15:0] b_30;
  wire [15:0] a_31;
  wire [15:0] b_31;
  wire [15:0] a_32;
  wire [15:0] b_32;
  wire [15:0] a_33;
  wire [15:0] b_33;
  wire [15:0] a_34;
  wire [15:0] b_34;
  wire [15:0] a_35;
  wire [15:0] b_35;
  wire [15:0] a_36;
  wire [15:0] b_36;
  wire [15:0] a_37;
  wire [15:0] b_37;
  wire [15:0] a_38;
  wire [15:0] b_38;
  wire [15:0] a_39;
  wire [15:0] b_39;
  wire [15:0] a_40;
  wire [15:0] b_40;
  wire [15:0] a_41;
  wire [15:0] b_41;
  wire [15:0] a_42;
  wire [15:0] b_42;
  wire [15:0] a_43;
  wire [15:0] b_43;
  wire [15:0] a_44;
  wire [15:0] b_44;
  wire [15:0] a_45;
  wire [15:0] b_45;
  wire [15:0] a_46;
  wire [15:0] b_46;
  wire [15:0] a_47;
  wire [15:0] b_47;
  wire [15:0] a_48;
  wire [15:0] b_48;
  wire [15:0] a_49;
  wire [15:0] b_49;
  wire [15:0] a_50;
  wire [15:0] b_50;
  wire [15:0] a_51;
  wire [15:0] b_51;
  wire [15:0] a_52;
  wire [15:0] b_52;
  wire [15:0] a_53;
  wire [15:0] b_53;
  wire [15:0] a_54;
  wire [15:0] b_54;
  wire [15:0] a_55;
  wire [15:0] b_55;
  wire [15:0] a_56;
  wire [15:0] b_56;
  wire [15:0] a_57;
  wire [15:0] b_57;
  wire [15:0] a_58;
  wire [15:0] b_58;
  wire [15:0] a_59;
  wire [15:0] b_59;
  wire [15:0] a_60;
  wire [15:0] b_60;
  wire [15:0] a_61;
  wire [15:0] b_61;
  wire [15:0] a_62;
  wire [15:0] b_62;
  wire [15:0] a_63;
  wire [15:0] b_63;
  wire [15:0] a_64;
  wire [15:0] b_64;
  wire [15:0] a_65;
  wire [15:0] b_65;
  wire [15:0] a_66;
  wire [15:0] b_66;
  wire [15:0] a_67;
  wire [15:0] b_67;
  wire [15:0] a_68;
  wire [15:0] b_68;
  wire [15:0] a_69;
  wire [15:0] b_69;
  wire [15:0] a_70;
  wire [15:0] b_70;
  wire [15:0] a_71;
  wire [15:0] b_71;
  wire [15:0] a_72;
  wire [15:0] b_72;
  wire [15:0] a_73;
  wire [15:0] b_73;
  wire [15:0] a_74;
  wire [15:0] b_74;
  wire [15:0] a_75;
  wire [15:0] b_75;
  wire [15:0] a_76;
  wire [15:0] b_76;
  wire [15:0] a_77;
  wire [15:0] b_77;
  wire [15:0] a_78;
  wire [15:0] b_78;
  wire [15:0] a_79;
  wire [15:0] b_79;
  wire [15:0] a_80;
  wire [15:0] b_80;
  wire [15:0] a_81;
  wire [15:0] b_81;
  wire [15:0] a_82;
  wire [15:0] b_82;
  wire [15:0] a_83;
  wire [15:0] b_83;
  reg [31:0] sum;
  reg [31:0] _RAND_0;
  reg [6:0] i;
  reg [31:0] _RAND_1;
  wire  _T_171;
  wire  _T_172;
  wire [15:0] _GEN_1;
  wire [15:0] _GEN_2;
  wire [15:0] _GEN_3;
  wire [15:0] _GEN_4;
  wire [15:0] _GEN_5;
  wire [15:0] _GEN_6;
  wire [15:0] _GEN_7;
  wire [15:0] _GEN_8;
  wire [15:0] _GEN_9;
  wire [15:0] _GEN_10;
  wire [15:0] _GEN_11;
  wire [15:0] _GEN_12;
  wire [15:0] _GEN_13;
  wire [15:0] _GEN_14;
  wire [15:0] _GEN_15;
  wire [15:0] _GEN_16;
  wire [15:0] _GEN_17;
  wire [15:0] _GEN_18;
  wire [15:0] _GEN_19;
  wire [15:0] _GEN_20;
  wire [15:0] _GEN_21;
  wire [15:0] _GEN_22;
  wire [15:0] _GEN_23;
  wire [15:0] _GEN_24;
  wire [15:0] _GEN_25;
  wire [15:0] _GEN_26;
  wire [15:0] _GEN_27;
  wire [15:0] _GEN_28;
  wire [15:0] _GEN_29;
  wire [15:0] _GEN_30;
  wire [15:0] _GEN_31;
  wire [15:0] _GEN_32;
  wire [15:0] _GEN_33;
  wire [15:0] _GEN_34;
  wire [15:0] _GEN_35;
  wire [15:0] _GEN_36;
  wire [15:0] _GEN_37;
  wire [15:0] _GEN_38;
  wire [15:0] _GEN_39;
  wire [15:0] _GEN_40;
  wire [15:0] _GEN_41;
  wire [15:0] _GEN_42;
  wire [15:0] _GEN_43;
  wire [15:0] _GEN_44;
  wire [15:0] _GEN_45;
  wire [15:0] _GEN_46;
  wire [15:0] _GEN_47;
  wire [15:0] _GEN_48;
  wire [15:0] _GEN_49;
  wire [15:0] _GEN_50;
  wire [15:0] _GEN_51;
  wire [15:0] _GEN_52;
  wire [15:0] _GEN_53;
  wire [15:0] _GEN_54;
  wire [15:0] _GEN_55;
  wire [15:0] _GEN_56;
  wire [15:0] _GEN_57;
  wire [15:0] _GEN_58;
  wire [15:0] _GEN_59;
  wire [15:0] _GEN_60;
  wire [15:0] _GEN_61;
  wire [15:0] _GEN_62;
  wire [15:0] _GEN_63;
  wire [15:0] _GEN_64;
  wire [15:0] _GEN_65;
  wire [15:0] _GEN_66;
  wire [15:0] _GEN_67;
  wire [15:0] _GEN_68;
  wire [15:0] _GEN_69;
  wire [15:0] _GEN_70;
  wire [15:0] _GEN_71;
  wire [15:0] _GEN_72;
  wire [15:0] _GEN_73;
  wire [15:0] _GEN_74;
  wire [15:0] _GEN_75;
  wire [15:0] _GEN_76;
  wire [15:0] _GEN_77;
  wire [15:0] _GEN_78;
  wire [15:0] _GEN_79;
  wire [15:0] _GEN_80;
  wire [15:0] _GEN_81;
  wire [15:0] _GEN_82;
  wire [15:0] _GEN_83;
  wire [15:0] _GEN_85;
  wire [15:0] _GEN_86;
  wire [15:0] _GEN_87;
  wire [15:0] _GEN_88;
  wire [15:0] _GEN_89;
  wire [15:0] _GEN_90;
  wire [15:0] _GEN_91;
  wire [15:0] _GEN_92;
  wire [15:0] _GEN_93;
  wire [15:0] _GEN_94;
  wire [15:0] _GEN_95;
  wire [15:0] _GEN_96;
  wire [15:0] _GEN_97;
  wire [15:0] _GEN_98;
  wire [15:0] _GEN_99;
  wire [15:0] _GEN_100;
  wire [15:0] _GEN_101;
  wire [15:0] _GEN_102;
  wire [15:0] _GEN_103;
  wire [15:0] _GEN_104;
  wire [15:0] _GEN_105;
  wire [15:0] _GEN_106;
  wire [15:0] _GEN_107;
  wire [15:0] _GEN_108;
  wire [15:0] _GEN_109;
  wire [15:0] _GEN_110;
  wire [15:0] _GEN_111;
  wire [15:0] _GEN_112;
  wire [15:0] _GEN_113;
  wire [15:0] _GEN_114;
  wire [15:0] _GEN_115;
  wire [15:0] _GEN_116;
  wire [15:0] _GEN_117;
  wire [15:0] _GEN_118;
  wire [15:0] _GEN_119;
  wire [15:0] _GEN_120;
  wire [15:0] _GEN_121;
  wire [15:0] _GEN_122;
  wire [15:0] _GEN_123;
  wire [15:0] _GEN_124;
  wire [15:0] _GEN_125;
  wire [15:0] _GEN_126;
  wire [15:0] _GEN_127;
  wire [15:0] _GEN_128;
  wire [15:0] _GEN_129;
  wire [15:0] _GEN_130;
  wire [15:0] _GEN_131;
  wire [15:0] _GEN_132;
  wire [15:0] _GEN_133;
  wire [15:0] _GEN_134;
  wire [15:0] _GEN_135;
  wire [15:0] _GEN_136;
  wire [15:0] _GEN_137;
  wire [15:0] _GEN_138;
  wire [15:0] _GEN_139;
  wire [15:0] _GEN_140;
  wire [15:0] _GEN_141;
  wire [15:0] _GEN_142;
  wire [15:0] _GEN_143;
  wire [15:0] _GEN_144;
  wire [15:0] _GEN_145;
  wire [15:0] _GEN_146;
  wire [15:0] _GEN_147;
  wire [15:0] _GEN_148;
  wire [15:0] _GEN_149;
  wire [15:0] _GEN_150;
  wire [15:0] _GEN_151;
  wire [15:0] _GEN_152;
  wire [15:0] _GEN_153;
  wire [15:0] _GEN_154;
  wire [15:0] _GEN_155;
  wire [15:0] _GEN_156;
  wire [15:0] _GEN_157;
  wire [15:0] _GEN_158;
  wire [15:0] _GEN_159;
  wire [15:0] _GEN_160;
  wire [15:0] _GEN_161;
  wire [15:0] _GEN_162;
  wire [15:0] _GEN_163;
  wire [15:0] _GEN_164;
  wire [15:0] _GEN_165;
  wire [15:0] _GEN_166;
  wire [15:0] _GEN_167;
  wire [31:0] _T_168;
  wire [32:0] _T_169;
  wire [7:0] _T_170;
  wire [7:0] _GEN_168;
  wire [32:0] _GEN_169;
  wire [7:0] _GEN_170;
  wire [31:0] _GEN_172;
  wire [32:0] _GEN_173;
  wire [32:0] _GEN_174;
  wire [7:0] _GEN_175;
  assign a_0 = io_a[15:0];
  assign b_0 = io_b[15:0];
  assign a_1 = io_a[31:16];
  assign b_1 = io_b[31:16];
  assign a_2 = io_a[47:32];
  assign b_2 = io_b[47:32];
  assign a_3 = io_a[63:48];
  assign b_3 = io_b[63:48];
  assign a_4 = io_a[79:64];
  assign b_4 = io_b[79:64];
  assign a_5 = io_a[95:80];
  assign b_5 = io_b[95:80];
  assign a_6 = io_a[111:96];
  assign b_6 = io_b[111:96];
  assign a_7 = io_a[127:112];
  assign b_7 = io_b[127:112];
  assign a_8 = io_a[143:128];
  assign b_8 = io_b[143:128];
  assign a_9 = io_a[159:144];
  assign b_9 = io_b[159:144];
  assign a_10 = io_a[175:160];
  assign b_10 = io_b[175:160];
  assign a_11 = io_a[191:176];
  assign b_11 = io_b[191:176];
  assign a_12 = io_a[207:192];
  assign b_12 = io_b[207:192];
  assign a_13 = io_a[223:208];
  assign b_13 = io_b[223:208];
  assign a_14 = io_a[239:224];
  assign b_14 = io_b[239:224];
  assign a_15 = io_a[255:240];
  assign b_15 = io_b[255:240];
  assign a_16 = io_a[271:256];
  assign b_16 = io_b[271:256];
  assign a_17 = io_a[287:272];
  assign b_17 = io_b[287:272];
  assign a_18 = io_a[303:288];
  assign b_18 = io_b[303:288];
  assign a_19 = io_a[319:304];
  assign b_19 = io_b[319:304];
  assign a_20 = io_a[335:320];
  assign b_20 = io_b[335:320];
  assign a_21 = io_a[351:336];
  assign b_21 = io_b[351:336];
  assign a_22 = io_a[367:352];
  assign b_22 = io_b[367:352];
  assign a_23 = io_a[383:368];
  assign b_23 = io_b[383:368];
  assign a_24 = io_a[399:384];
  assign b_24 = io_b[399:384];
  assign a_25 = io_a[415:400];
  assign b_25 = io_b[415:400];
  assign a_26 = io_a[431:416];
  assign b_26 = io_b[431:416];
  assign a_27 = io_a[447:432];
  assign b_27 = io_b[447:432];
  assign a_28 = io_a[463:448];
  assign b_28 = io_b[463:448];
  assign a_29 = io_a[479:464];
  assign b_29 = io_b[479:464];
  assign a_30 = io_a[495:480];
  assign b_30 = io_b[495:480];
  assign a_31 = io_a[511:496];
  assign b_31 = io_b[511:496];
  assign a_32 = io_a[527:512];
  assign b_32 = io_b[527:512];
  assign a_33 = io_a[543:528];
  assign b_33 = io_b[543:528];
  assign a_34 = io_a[559:544];
  assign b_34 = io_b[559:544];
  assign a_35 = io_a[575:560];
  assign b_35 = io_b[575:560];
  assign a_36 = io_a[591:576];
  assign b_36 = io_b[591:576];
  assign a_37 = io_a[607:592];
  assign b_37 = io_b[607:592];
  assign a_38 = io_a[623:608];
  assign b_38 = io_b[623:608];
  assign a_39 = io_a[639:624];
  assign b_39 = io_b[639:624];
  assign a_40 = io_a[655:640];
  assign b_40 = io_b[655:640];
  assign a_41 = io_a[671:656];
  assign b_41 = io_b[671:656];
  assign a_42 = io_a[687:672];
  assign b_42 = io_b[687:672];
  assign a_43 = io_a[703:688];
  assign b_43 = io_b[703:688];
  assign a_44 = io_a[719:704];
  assign b_44 = io_b[719:704];
  assign a_45 = io_a[735:720];
  assign b_45 = io_b[735:720];
  assign a_46 = io_a[751:736];
  assign b_46 = io_b[751:736];
  assign a_47 = io_a[767:752];
  assign b_47 = io_b[767:752];
  assign a_48 = io_a[783:768];
  assign b_48 = io_b[783:768];
  assign a_49 = io_a[799:784];
  assign b_49 = io_b[799:784];
  assign a_50 = io_a[815:800];
  assign b_50 = io_b[815:800];
  assign a_51 = io_a[831:816];
  assign b_51 = io_b[831:816];
  assign a_52 = io_a[847:832];
  assign b_52 = io_b[847:832];
  assign a_53 = io_a[863:848];
  assign b_53 = io_b[863:848];
  assign a_54 = io_a[879:864];
  assign b_54 = io_b[879:864];
  assign a_55 = io_a[895:880];
  assign b_55 = io_b[895:880];
  assign a_56 = io_a[911:896];
  assign b_56 = io_b[911:896];
  assign a_57 = io_a[927:912];
  assign b_57 = io_b[927:912];
  assign a_58 = io_a[943:928];
  assign b_58 = io_b[943:928];
  assign a_59 = io_a[959:944];
  assign b_59 = io_b[959:944];
  assign a_60 = io_a[975:960];
  assign b_60 = io_b[975:960];
  assign a_61 = io_a[991:976];
  assign b_61 = io_b[991:976];
  assign a_62 = io_a[1007:992];
  assign b_62 = io_b[1007:992];
  assign a_63 = io_a[1023:1008];
  assign b_63 = io_b[1023:1008];
  assign a_64 = io_a[1039:1024];
  assign b_64 = io_b[1039:1024];
  assign a_65 = io_a[1055:1040];
  assign b_65 = io_b[1055:1040];
  assign a_66 = io_a[1071:1056];
  assign b_66 = io_b[1071:1056];
  assign a_67 = io_a[1087:1072];
  assign b_67 = io_b[1087:1072];
  assign a_68 = io_a[1103:1088];
  assign b_68 = io_b[1103:1088];
  assign a_69 = io_a[1119:1104];
  assign b_69 = io_b[1119:1104];
  assign a_70 = io_a[1135:1120];
  assign b_70 = io_b[1135:1120];
  assign a_71 = io_a[1151:1136];
  assign b_71 = io_b[1151:1136];
  assign a_72 = io_a[1167:1152];
  assign b_72 = io_b[1167:1152];
  assign a_73 = io_a[1183:1168];
  assign b_73 = io_b[1183:1168];
  assign a_74 = io_a[1199:1184];
  assign b_74 = io_b[1199:1184];
  assign a_75 = io_a[1215:1200];
  assign b_75 = io_b[1215:1200];
  assign a_76 = io_a[1231:1216];
  assign b_76 = io_b[1231:1216];
  assign a_77 = io_a[1247:1232];
  assign b_77 = io_b[1247:1232];
  assign a_78 = io_a[1263:1248];
  assign b_78 = io_b[1263:1248];
  assign a_79 = io_a[1279:1264];
  assign b_79 = io_b[1279:1264];
  assign a_80 = io_a[1295:1280];
  assign b_80 = io_b[1295:1280];
  assign a_81 = io_a[1311:1296];
  assign b_81 = io_b[1311:1296];
  assign a_82 = io_a[1327:1312];
  assign b_82 = io_b[1327:1312];
  assign a_83 = io_a[1343:1328];
  assign b_83 = io_b[1343:1328];
  assign _T_171 = i == 7'h54;
  assign _T_172 = i != 7'h0;
  assign _GEN_1 = 7'h1 == i ? a_1 : a_0;
  assign _GEN_2 = 7'h2 == i ? a_2 : _GEN_1;
  assign _GEN_3 = 7'h3 == i ? a_3 : _GEN_2;
  assign _GEN_4 = 7'h4 == i ? a_4 : _GEN_3;
  assign _GEN_5 = 7'h5 == i ? a_5 : _GEN_4;
  assign _GEN_6 = 7'h6 == i ? a_6 : _GEN_5;
  assign _GEN_7 = 7'h7 == i ? a_7 : _GEN_6;
  assign _GEN_8 = 7'h8 == i ? a_8 : _GEN_7;
  assign _GEN_9 = 7'h9 == i ? a_9 : _GEN_8;
  assign _GEN_10 = 7'ha == i ? a_10 : _GEN_9;
  assign _GEN_11 = 7'hb == i ? a_11 : _GEN_10;
  assign _GEN_12 = 7'hc == i ? a_12 : _GEN_11;
  assign _GEN_13 = 7'hd == i ? a_13 : _GEN_12;
  assign _GEN_14 = 7'he == i ? a_14 : _GEN_13;
  assign _GEN_15 = 7'hf == i ? a_15 : _GEN_14;
  assign _GEN_16 = 7'h10 == i ? a_16 : _GEN_15;
  assign _GEN_17 = 7'h11 == i ? a_17 : _GEN_16;
  assign _GEN_18 = 7'h12 == i ? a_18 : _GEN_17;
  assign _GEN_19 = 7'h13 == i ? a_19 : _GEN_18;
  assign _GEN_20 = 7'h14 == i ? a_20 : _GEN_19;
  assign _GEN_21 = 7'h15 == i ? a_21 : _GEN_20;
  assign _GEN_22 = 7'h16 == i ? a_22 : _GEN_21;
  assign _GEN_23 = 7'h17 == i ? a_23 : _GEN_22;
  assign _GEN_24 = 7'h18 == i ? a_24 : _GEN_23;
  assign _GEN_25 = 7'h19 == i ? a_25 : _GEN_24;
  assign _GEN_26 = 7'h1a == i ? a_26 : _GEN_25;
  assign _GEN_27 = 7'h1b == i ? a_27 : _GEN_26;
  assign _GEN_28 = 7'h1c == i ? a_28 : _GEN_27;
  assign _GEN_29 = 7'h1d == i ? a_29 : _GEN_28;
  assign _GEN_30 = 7'h1e == i ? a_30 : _GEN_29;
  assign _GEN_31 = 7'h1f == i ? a_31 : _GEN_30;
  assign _GEN_32 = 7'h20 == i ? a_32 : _GEN_31;
  assign _GEN_33 = 7'h21 == i ? a_33 : _GEN_32;
  assign _GEN_34 = 7'h22 == i ? a_34 : _GEN_33;
  assign _GEN_35 = 7'h23 == i ? a_35 : _GEN_34;
  assign _GEN_36 = 7'h24 == i ? a_36 : _GEN_35;
  assign _GEN_37 = 7'h25 == i ? a_37 : _GEN_36;
  assign _GEN_38 = 7'h26 == i ? a_38 : _GEN_37;
  assign _GEN_39 = 7'h27 == i ? a_39 : _GEN_38;
  assign _GEN_40 = 7'h28 == i ? a_40 : _GEN_39;
  assign _GEN_41 = 7'h29 == i ? a_41 : _GEN_40;
  assign _GEN_42 = 7'h2a == i ? a_42 : _GEN_41;
  assign _GEN_43 = 7'h2b == i ? a_43 : _GEN_42;
  assign _GEN_44 = 7'h2c == i ? a_44 : _GEN_43;
  assign _GEN_45 = 7'h2d == i ? a_45 : _GEN_44;
  assign _GEN_46 = 7'h2e == i ? a_46 : _GEN_45;
  assign _GEN_47 = 7'h2f == i ? a_47 : _GEN_46;
  assign _GEN_48 = 7'h30 == i ? a_48 : _GEN_47;
  assign _GEN_49 = 7'h31 == i ? a_49 : _GEN_48;
  assign _GEN_50 = 7'h32 == i ? a_50 : _GEN_49;
  assign _GEN_51 = 7'h33 == i ? a_51 : _GEN_50;
  assign _GEN_52 = 7'h34 == i ? a_52 : _GEN_51;
  assign _GEN_53 = 7'h35 == i ? a_53 : _GEN_52;
  assign _GEN_54 = 7'h36 == i ? a_54 : _GEN_53;
  assign _GEN_55 = 7'h37 == i ? a_55 : _GEN_54;
  assign _GEN_56 = 7'h38 == i ? a_56 : _GEN_55;
  assign _GEN_57 = 7'h39 == i ? a_57 : _GEN_56;
  assign _GEN_58 = 7'h3a == i ? a_58 : _GEN_57;
  assign _GEN_59 = 7'h3b == i ? a_59 : _GEN_58;
  assign _GEN_60 = 7'h3c == i ? a_60 : _GEN_59;
  assign _GEN_61 = 7'h3d == i ? a_61 : _GEN_60;
  assign _GEN_62 = 7'h3e == i ? a_62 : _GEN_61;
  assign _GEN_63 = 7'h3f == i ? a_63 : _GEN_62;
  assign _GEN_64 = 7'h40 == i ? a_64 : _GEN_63;
  assign _GEN_65 = 7'h41 == i ? a_65 : _GEN_64;
  assign _GEN_66 = 7'h42 == i ? a_66 : _GEN_65;
  assign _GEN_67 = 7'h43 == i ? a_67 : _GEN_66;
  assign _GEN_68 = 7'h44 == i ? a_68 : _GEN_67;
  assign _GEN_69 = 7'h45 == i ? a_69 : _GEN_68;
  assign _GEN_70 = 7'h46 == i ? a_70 : _GEN_69;
  assign _GEN_71 = 7'h47 == i ? a_71 : _GEN_70;
  assign _GEN_72 = 7'h48 == i ? a_72 : _GEN_71;
  assign _GEN_73 = 7'h49 == i ? a_73 : _GEN_72;
  assign _GEN_74 = 7'h4a == i ? a_74 : _GEN_73;
  assign _GEN_75 = 7'h4b == i ? a_75 : _GEN_74;
  assign _GEN_76 = 7'h4c == i ? a_76 : _GEN_75;
  assign _GEN_77 = 7'h4d == i ? a_77 : _GEN_76;
  assign _GEN_78 = 7'h4e == i ? a_78 : _GEN_77;
  assign _GEN_79 = 7'h4f == i ? a_79 : _GEN_78;
  assign _GEN_80 = 7'h50 == i ? a_80 : _GEN_79;
  assign _GEN_81 = 7'h51 == i ? a_81 : _GEN_80;
  assign _GEN_82 = 7'h52 == i ? a_82 : _GEN_81;
  assign _GEN_83 = 7'h53 == i ? a_83 : _GEN_82;
  assign _GEN_85 = 7'h1 == i ? b_1 : b_0;
  assign _GEN_86 = 7'h2 == i ? b_2 : _GEN_85;
  assign _GEN_87 = 7'h3 == i ? b_3 : _GEN_86;
  assign _GEN_88 = 7'h4 == i ? b_4 : _GEN_87;
  assign _GEN_89 = 7'h5 == i ? b_5 : _GEN_88;
  assign _GEN_90 = 7'h6 == i ? b_6 : _GEN_89;
  assign _GEN_91 = 7'h7 == i ? b_7 : _GEN_90;
  assign _GEN_92 = 7'h8 == i ? b_8 : _GEN_91;
  assign _GEN_93 = 7'h9 == i ? b_9 : _GEN_92;
  assign _GEN_94 = 7'ha == i ? b_10 : _GEN_93;
  assign _GEN_95 = 7'hb == i ? b_11 : _GEN_94;
  assign _GEN_96 = 7'hc == i ? b_12 : _GEN_95;
  assign _GEN_97 = 7'hd == i ? b_13 : _GEN_96;
  assign _GEN_98 = 7'he == i ? b_14 : _GEN_97;
  assign _GEN_99 = 7'hf == i ? b_15 : _GEN_98;
  assign _GEN_100 = 7'h10 == i ? b_16 : _GEN_99;
  assign _GEN_101 = 7'h11 == i ? b_17 : _GEN_100;
  assign _GEN_102 = 7'h12 == i ? b_18 : _GEN_101;
  assign _GEN_103 = 7'h13 == i ? b_19 : _GEN_102;
  assign _GEN_104 = 7'h14 == i ? b_20 : _GEN_103;
  assign _GEN_105 = 7'h15 == i ? b_21 : _GEN_104;
  assign _GEN_106 = 7'h16 == i ? b_22 : _GEN_105;
  assign _GEN_107 = 7'h17 == i ? b_23 : _GEN_106;
  assign _GEN_108 = 7'h18 == i ? b_24 : _GEN_107;
  assign _GEN_109 = 7'h19 == i ? b_25 : _GEN_108;
  assign _GEN_110 = 7'h1a == i ? b_26 : _GEN_109;
  assign _GEN_111 = 7'h1b == i ? b_27 : _GEN_110;
  assign _GEN_112 = 7'h1c == i ? b_28 : _GEN_111;
  assign _GEN_113 = 7'h1d == i ? b_29 : _GEN_112;
  assign _GEN_114 = 7'h1e == i ? b_30 : _GEN_113;
  assign _GEN_115 = 7'h1f == i ? b_31 : _GEN_114;
  assign _GEN_116 = 7'h20 == i ? b_32 : _GEN_115;
  assign _GEN_117 = 7'h21 == i ? b_33 : _GEN_116;
  assign _GEN_118 = 7'h22 == i ? b_34 : _GEN_117;
  assign _GEN_119 = 7'h23 == i ? b_35 : _GEN_118;
  assign _GEN_120 = 7'h24 == i ? b_36 : _GEN_119;
  assign _GEN_121 = 7'h25 == i ? b_37 : _GEN_120;
  assign _GEN_122 = 7'h26 == i ? b_38 : _GEN_121;
  assign _GEN_123 = 7'h27 == i ? b_39 : _GEN_122;
  assign _GEN_124 = 7'h28 == i ? b_40 : _GEN_123;
  assign _GEN_125 = 7'h29 == i ? b_41 : _GEN_124;
  assign _GEN_126 = 7'h2a == i ? b_42 : _GEN_125;
  assign _GEN_127 = 7'h2b == i ? b_43 : _GEN_126;
  assign _GEN_128 = 7'h2c == i ? b_44 : _GEN_127;
  assign _GEN_129 = 7'h2d == i ? b_45 : _GEN_128;
  assign _GEN_130 = 7'h2e == i ? b_46 : _GEN_129;
  assign _GEN_131 = 7'h2f == i ? b_47 : _GEN_130;
  assign _GEN_132 = 7'h30 == i ? b_48 : _GEN_131;
  assign _GEN_133 = 7'h31 == i ? b_49 : _GEN_132;
  assign _GEN_134 = 7'h32 == i ? b_50 : _GEN_133;
  assign _GEN_135 = 7'h33 == i ? b_51 : _GEN_134;
  assign _GEN_136 = 7'h34 == i ? b_52 : _GEN_135;
  assign _GEN_137 = 7'h35 == i ? b_53 : _GEN_136;
  assign _GEN_138 = 7'h36 == i ? b_54 : _GEN_137;
  assign _GEN_139 = 7'h37 == i ? b_55 : _GEN_138;
  assign _GEN_140 = 7'h38 == i ? b_56 : _GEN_139;
  assign _GEN_141 = 7'h39 == i ? b_57 : _GEN_140;
  assign _GEN_142 = 7'h3a == i ? b_58 : _GEN_141;
  assign _GEN_143 = 7'h3b == i ? b_59 : _GEN_142;
  assign _GEN_144 = 7'h3c == i ? b_60 : _GEN_143;
  assign _GEN_145 = 7'h3d == i ? b_61 : _GEN_144;
  assign _GEN_146 = 7'h3e == i ? b_62 : _GEN_145;
  assign _GEN_147 = 7'h3f == i ? b_63 : _GEN_146;
  assign _GEN_148 = 7'h40 == i ? b_64 : _GEN_147;
  assign _GEN_149 = 7'h41 == i ? b_65 : _GEN_148;
  assign _GEN_150 = 7'h42 == i ? b_66 : _GEN_149;
  assign _GEN_151 = 7'h43 == i ? b_67 : _GEN_150;
  assign _GEN_152 = 7'h44 == i ? b_68 : _GEN_151;
  assign _GEN_153 = 7'h45 == i ? b_69 : _GEN_152;
  assign _GEN_154 = 7'h46 == i ? b_70 : _GEN_153;
  assign _GEN_155 = 7'h47 == i ? b_71 : _GEN_154;
  assign _GEN_156 = 7'h48 == i ? b_72 : _GEN_155;
  assign _GEN_157 = 7'h49 == i ? b_73 : _GEN_156;
  assign _GEN_158 = 7'h4a == i ? b_74 : _GEN_157;
  assign _GEN_159 = 7'h4b == i ? b_75 : _GEN_158;
  assign _GEN_160 = 7'h4c == i ? b_76 : _GEN_159;
  assign _GEN_161 = 7'h4d == i ? b_77 : _GEN_160;
  assign _GEN_162 = 7'h4e == i ? b_78 : _GEN_161;
  assign _GEN_163 = 7'h4f == i ? b_79 : _GEN_162;
  assign _GEN_164 = 7'h50 == i ? b_80 : _GEN_163;
  assign _GEN_165 = 7'h51 == i ? b_81 : _GEN_164;
  assign _GEN_166 = 7'h52 == i ? b_82 : _GEN_165;
  assign _GEN_167 = 7'h53 == i ? b_83 : _GEN_166;
  assign _T_168 = _GEN_83 * _GEN_167;
  assign _T_169 = sum + _T_168;
  assign _T_170 = i + 7'h1;
  assign _GEN_168 = _T_172 ? _T_170 : 8'h0;
  assign _GEN_169 = _T_172 ? _T_169 : 33'h0;
  assign _GEN_170 = _T_171 ? 8'h0 : _GEN_168;
  assign _GEN_172 = _T_171 ? sum : 32'h0;
  assign _GEN_173 = _T_171 ? 33'h0 : _GEN_169;
  assign _GEN_174 = io_rdy ? _T_169 : _GEN_173;
  assign _GEN_175 = io_rdy ? _T_170 : _GEN_170;
  assign io_q = io_rdy ? 32'h0 : _GEN_172;
  assign io_v = io_rdy ? 1'h0 : _T_171;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sum = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  i = _RAND_1[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      sum <= 32'h0;
    end else begin
      sum <= _GEN_174[31:0];
    end
    if (reset) begin
      i <= 7'h0;
    end else begin
      i <= _GEN_175[6:0];
    end
  end
endmodule
module Node_104(
  input           clock,
  input           reset,
  input  [1343:0] io_d_in,
  input  [1343:0] io_w,
  input           io_rdy,
  input  [15:0]   io_bias,
  output [15:0]   io_d_out,
  output          io_v
);
  wire  muladdc_clock;
  wire  muladdc_reset;
  wire [1343:0] muladdc_io_a;
  wire [1343:0] muladdc_io_b;
  wire  muladdc_io_rdy;
  wire [31:0] muladdc_io_q;
  wire  muladdc_io_v;
  wire [31:0] act_io_q;
  wire [15:0] act_io_bias;
  wire  act_io_v_in;
  wire [15:0] act_io_d;
  wire  act_io_v_out;
  Mac_104 muladdc (
    .clock(muladdc_clock),
    .reset(muladdc_reset),
    .io_a(muladdc_io_a),
    .io_b(muladdc_io_b),
    .io_rdy(muladdc_io_rdy),
    .io_q(muladdc_io_q),
    .io_v(muladdc_io_v)
  );
  ReLU act (
    .io_q(act_io_q),
    .io_bias(act_io_bias),
    .io_v_in(act_io_v_in),
    .io_d(act_io_d),
    .io_v_out(act_io_v_out)
  );
  assign io_d_out = act_io_d;
  assign io_v = act_io_v_out;
  assign muladdc_clock = clock;
  assign muladdc_reset = reset;
  assign muladdc_io_a = io_d_in;
  assign muladdc_io_b = io_w;
  assign muladdc_io_rdy = io_rdy;
  assign act_io_q = muladdc_io_q;
  assign act_io_bias = io_bias;
  assign act_io_v_in = muladdc_io_v;
endmodule
module FC3(
  input           clock,
  input           reset,
  input  [15:0]   io_d_in,
  input  [1343:0] io_w_in,
  input  [159:0]  io_bias,
  input           io_rdy,
  input           io_done,
  output [15:0]   io_d_out,
  output          io_v,
  output          io_fc2_done
);
  wire  in_channel_clock;
  wire  in_channel_reset;
  wire [15:0] in_channel_io_d_in;
  wire  in_channel_io_en;
  wire [1343:0] in_channel_io_d_out;
  wire  conv_node3_clock;
  wire  conv_node3_reset;
  wire [1343:0] conv_node3_io_d_in;
  wire [1343:0] conv_node3_io_w;
  wire  conv_node3_io_rdy;
  wire [15:0] conv_node3_io_bias;
  wire [15:0] conv_node3_io_d_out;
  wire  conv_node3_io_v;
  reg  rdy;
  reg [31:0] _RAND_0;
  reg [1343:0] store;
  reg [1343:0] _RAND_1;
  reg  first_rdy;
  reg [31:0] _RAND_2;
  reg [15:0] in_counter;
  reg [31:0] _RAND_3;
  wire  _T;
  wire [16:0] _T_1;
  wire [16:0] _GEN_0;
  wire [16:0] _GEN_1;
  reg  is_done;
  reg [31:0] _RAND_4;
  wire  _GEN_4;
  wire  _T_2;
  ShiftRegister_23 in_channel (
    .clock(in_channel_clock),
    .reset(in_channel_reset),
    .io_d_in(in_channel_io_d_in),
    .io_en(in_channel_io_en),
    .io_d_out(in_channel_io_d_out)
  );
  Node_104 conv_node3 (
    .clock(conv_node3_clock),
    .reset(conv_node3_reset),
    .io_d_in(conv_node3_io_d_in),
    .io_w(conv_node3_io_w),
    .io_rdy(conv_node3_io_rdy),
    .io_bias(conv_node3_io_bias),
    .io_d_out(conv_node3_io_d_out),
    .io_v(conv_node3_io_v)
  );
  assign _T = in_counter == 16'h54;
  assign _T_1 = in_counter + 16'h1;
  assign _GEN_0 = io_rdy ? _T_1 : {{1'd0}, in_counter};
  assign _GEN_1 = _T ? 17'h0 : _GEN_0;
  assign _GEN_4 = io_done | is_done;
  assign _T_2 = first_rdy | conv_node3_io_v;
  assign io_d_out = conv_node3_io_d_out;
  assign io_v = conv_node3_io_v;
  assign io_fc2_done = in_counter == 16'h54;
  assign in_channel_clock = clock;
  assign in_channel_reset = reset;
  assign in_channel_io_d_in = io_d_in;
  assign in_channel_io_en = io_rdy;
  assign conv_node3_clock = clock;
  assign conv_node3_reset = reset;
  assign conv_node3_io_d_in = store;
  assign conv_node3_io_w = io_w_in;
  assign conv_node3_io_rdy = rdy;
  assign conv_node3_io_bias = io_bias[15:0];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rdy = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {42{`RANDOM}};
  store = _RAND_1[1343:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  first_rdy = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_counter = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  is_done = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      rdy <= 1'h0;
    end else if (is_done) begin
      rdy <= 1'h0;
    end else begin
      rdy <= _T_2;
    end
    if (reset) begin
      store <= 1344'h0;
    end else if (_T) begin
      store <= in_channel_io_d_out;
    end
    if (reset) begin
      first_rdy <= 1'h0;
    end else begin
      first_rdy <= _T;
    end
    if (reset) begin
      in_counter <= 16'h0;
    end else begin
      in_counter <= _GEN_1[15:0];
    end
    if (reset) begin
      is_done <= 1'h0;
    end else begin
      is_done <= _GEN_4;
    end
  end
endmodule
module Top(
  input           clock,
  input           reset,
  input  [399:0]  io_d_in,
  input  [399:0]  io_w_in_0,
  input  [399:0]  io_w_in_1,
  input  [399:0]  io_w_in_2,
  input  [399:0]  io_w_in_3,
  input  [399:0]  io_w_in_4,
  input  [399:0]  io_w_in_5,
  input  [95:0]   io_bias,
  input           io_rdy,
  output          io_v,
  output          io_c3_v,
  output          io_pool_v,
  input  [3199:0] io_fc1_wa_in,
  input  [3199:0] io_fc1_wb_in,
  input  [15:0]   io_fc1_bias,
  input           io_fc1_rom_rdy,
  output          io_fc1_v,
  output          io_fc1_fc_v,
  input  [1919:0] io_fc2_w_in,
  input  [15:0]   io_fc2_bias,
  input           io_fc2_rom_rdy,
  output          io_fc2_v,
  output          io_fc2_fc_v,
  input  [1343:0] io_fc3_w_in,
  input  [15:0]   io_fc3_bias,
  input           io_fc3_rom_rdy,
  output [15:0]   io_fc3_d_out,
  output          io_fc3_v,
  output          io_fc3_fc_v
);
  wire  t1_clock;
  wire  t1_reset;
  wire [399:0] t1_io_d_in;
  wire [399:0] t1_io_w_in_0;
  wire [399:0] t1_io_w_in_1;
  wire [399:0] t1_io_w_in_2;
  wire [399:0] t1_io_w_in_3;
  wire [399:0] t1_io_w_in_4;
  wire [399:0] t1_io_w_in_5;
  wire [95:0] t1_io_bias;
  wire  t1_io_rdy;
  wire  t1_io_v;
  wire [15:0] t1_io_d_out_0;
  wire [15:0] t1_io_d_out_1;
  wire [15:0] t1_io_d_out_2;
  wire [15:0] t1_io_d_out_3;
  wire [15:0] t1_io_d_out_4;
  wire [15:0] t1_io_d_out_5;
  wire  t1_io_pool_v;
  wire  t2_clock;
  wire  t2_reset;
  wire [15:0] t2_io_d_in_0;
  wire [15:0] t2_io_d_in_1;
  wire [15:0] t2_io_d_in_2;
  wire [15:0] t2_io_d_in_3;
  wire [15:0] t2_io_d_in_4;
  wire [15:0] t2_io_d_in_5;
  wire  t2_io_rdy;
  wire  t2_io_c3_v;
  wire [15:0] t2_io_d_out_0;
  wire [15:0] t2_io_d_out_1;
  wire [15:0] t2_io_d_out_2;
  wire [15:0] t2_io_d_out_3;
  wire [15:0] t2_io_d_out_4;
  wire [15:0] t2_io_d_out_5;
  wire [15:0] t2_io_d_out_6;
  wire [15:0] t2_io_d_out_7;
  wire [15:0] t2_io_d_out_8;
  wire [15:0] t2_io_d_out_9;
  wire [15:0] t2_io_d_out_10;
  wire [15:0] t2_io_d_out_11;
  wire [15:0] t2_io_d_out_12;
  wire [15:0] t2_io_d_out_13;
  wire [15:0] t2_io_d_out_14;
  wire [15:0] t2_io_d_out_15;
  wire  c2mp_clock;
  wire  c2mp_reset;
  wire [15:0] c2mp_io_d_in_0;
  wire [15:0] c2mp_io_d_in_1;
  wire [15:0] c2mp_io_d_in_2;
  wire [15:0] c2mp_io_d_in_3;
  wire [15:0] c2mp_io_d_in_4;
  wire [15:0] c2mp_io_d_in_5;
  wire [15:0] c2mp_io_d_in_6;
  wire [15:0] c2mp_io_d_in_7;
  wire [15:0] c2mp_io_d_in_8;
  wire [15:0] c2mp_io_d_in_9;
  wire [15:0] c2mp_io_d_in_10;
  wire [15:0] c2mp_io_d_in_11;
  wire [15:0] c2mp_io_d_in_12;
  wire [15:0] c2mp_io_d_in_13;
  wire [15:0] c2mp_io_d_in_14;
  wire [15:0] c2mp_io_d_in_15;
  wire  c2mp_io_rdy;
  wire [15:0] c2mp_io_d_out_0;
  wire [15:0] c2mp_io_d_out_1;
  wire [15:0] c2mp_io_d_out_2;
  wire [15:0] c2mp_io_d_out_3;
  wire [15:0] c2mp_io_d_out_4;
  wire [15:0] c2mp_io_d_out_5;
  wire [15:0] c2mp_io_d_out_6;
  wire [15:0] c2mp_io_d_out_7;
  wire [15:0] c2mp_io_d_out_8;
  wire [15:0] c2mp_io_d_out_9;
  wire [15:0] c2mp_io_d_out_10;
  wire [15:0] c2mp_io_d_out_11;
  wire [15:0] c2mp_io_d_out_12;
  wire [15:0] c2mp_io_d_out_13;
  wire [15:0] c2mp_io_d_out_14;
  wire [15:0] c2mp_io_d_out_15;
  wire  c2mp_io_pool_v;
  wire  f1_clock;
  wire  f1_reset;
  wire [15:0] f1_io_d_in_0;
  wire [15:0] f1_io_d_in_1;
  wire [15:0] f1_io_d_in_2;
  wire [15:0] f1_io_d_in_3;
  wire [15:0] f1_io_d_in_4;
  wire [15:0] f1_io_d_in_5;
  wire [15:0] f1_io_d_in_6;
  wire [15:0] f1_io_d_in_7;
  wire [15:0] f1_io_d_in_8;
  wire [15:0] f1_io_d_in_9;
  wire [15:0] f1_io_d_in_10;
  wire [15:0] f1_io_d_in_11;
  wire [15:0] f1_io_d_in_12;
  wire [15:0] f1_io_d_in_13;
  wire [15:0] f1_io_d_in_14;
  wire [15:0] f1_io_d_in_15;
  wire [3199:0] f1_io_wa_in;
  wire [3199:0] f1_io_wb_in;
  wire [15:0] f1_io_bias;
  wire  f1_io_rdy;
  wire  f1_io_done;
  wire [15:0] f1_io_d_out;
  wire  f1_io_v;
  wire  f2_clock;
  wire  f2_reset;
  wire [15:0] f2_io_d_in;
  wire [1919:0] f2_io_w_in;
  wire [15:0] f2_io_bias;
  wire  f2_io_rdy;
  wire  f2_io_done;
  wire [15:0] f2_io_d_out;
  wire  f2_io_v;
  wire  f2_io_fc1_done;
  wire  f3_clock;
  wire  f3_reset;
  wire [15:0] f3_io_d_in;
  wire [1343:0] f3_io_w_in;
  wire [159:0] f3_io_bias;
  wire  f3_io_rdy;
  wire  f3_io_done;
  wire [15:0] f3_io_d_out;
  wire  f3_io_v;
  wire  f3_io_fc2_done;
  reg  delay_c3;
  reg [31:0] _RAND_0;
  reg [15:0] fc3_counter;
  reg [31:0] _RAND_1;
  wire  _T;
  wire [16:0] _T_1;
  wire [16:0] _GEN_0;
  wire [16:0] _GEN_1;
  Tile t1 (
    .clock(t1_clock),
    .reset(t1_reset),
    .io_d_in(t1_io_d_in),
    .io_w_in_0(t1_io_w_in_0),
    .io_w_in_1(t1_io_w_in_1),
    .io_w_in_2(t1_io_w_in_2),
    .io_w_in_3(t1_io_w_in_3),
    .io_w_in_4(t1_io_w_in_4),
    .io_w_in_5(t1_io_w_in_5),
    .io_bias(t1_io_bias),
    .io_rdy(t1_io_rdy),
    .io_v(t1_io_v),
    .io_d_out_0(t1_io_d_out_0),
    .io_d_out_1(t1_io_d_out_1),
    .io_d_out_2(t1_io_d_out_2),
    .io_d_out_3(t1_io_d_out_3),
    .io_d_out_4(t1_io_d_out_4),
    .io_d_out_5(t1_io_d_out_5),
    .io_pool_v(t1_io_pool_v)
  );
  Tile2 t2 (
    .clock(t2_clock),
    .reset(t2_reset),
    .io_d_in_0(t2_io_d_in_0),
    .io_d_in_1(t2_io_d_in_1),
    .io_d_in_2(t2_io_d_in_2),
    .io_d_in_3(t2_io_d_in_3),
    .io_d_in_4(t2_io_d_in_4),
    .io_d_in_5(t2_io_d_in_5),
    .io_rdy(t2_io_rdy),
    .io_c3_v(t2_io_c3_v),
    .io_d_out_0(t2_io_d_out_0),
    .io_d_out_1(t2_io_d_out_1),
    .io_d_out_2(t2_io_d_out_2),
    .io_d_out_3(t2_io_d_out_3),
    .io_d_out_4(t2_io_d_out_4),
    .io_d_out_5(t2_io_d_out_5),
    .io_d_out_6(t2_io_d_out_6),
    .io_d_out_7(t2_io_d_out_7),
    .io_d_out_8(t2_io_d_out_8),
    .io_d_out_9(t2_io_d_out_9),
    .io_d_out_10(t2_io_d_out_10),
    .io_d_out_11(t2_io_d_out_11),
    .io_d_out_12(t2_io_d_out_12),
    .io_d_out_13(t2_io_d_out_13),
    .io_d_out_14(t2_io_d_out_14),
    .io_d_out_15(t2_io_d_out_15)
  );
  C2MaxPool c2mp (
    .clock(c2mp_clock),
    .reset(c2mp_reset),
    .io_d_in_0(c2mp_io_d_in_0),
    .io_d_in_1(c2mp_io_d_in_1),
    .io_d_in_2(c2mp_io_d_in_2),
    .io_d_in_3(c2mp_io_d_in_3),
    .io_d_in_4(c2mp_io_d_in_4),
    .io_d_in_5(c2mp_io_d_in_5),
    .io_d_in_6(c2mp_io_d_in_6),
    .io_d_in_7(c2mp_io_d_in_7),
    .io_d_in_8(c2mp_io_d_in_8),
    .io_d_in_9(c2mp_io_d_in_9),
    .io_d_in_10(c2mp_io_d_in_10),
    .io_d_in_11(c2mp_io_d_in_11),
    .io_d_in_12(c2mp_io_d_in_12),
    .io_d_in_13(c2mp_io_d_in_13),
    .io_d_in_14(c2mp_io_d_in_14),
    .io_d_in_15(c2mp_io_d_in_15),
    .io_rdy(c2mp_io_rdy),
    .io_d_out_0(c2mp_io_d_out_0),
    .io_d_out_1(c2mp_io_d_out_1),
    .io_d_out_2(c2mp_io_d_out_2),
    .io_d_out_3(c2mp_io_d_out_3),
    .io_d_out_4(c2mp_io_d_out_4),
    .io_d_out_5(c2mp_io_d_out_5),
    .io_d_out_6(c2mp_io_d_out_6),
    .io_d_out_7(c2mp_io_d_out_7),
    .io_d_out_8(c2mp_io_d_out_8),
    .io_d_out_9(c2mp_io_d_out_9),
    .io_d_out_10(c2mp_io_d_out_10),
    .io_d_out_11(c2mp_io_d_out_11),
    .io_d_out_12(c2mp_io_d_out_12),
    .io_d_out_13(c2mp_io_d_out_13),
    .io_d_out_14(c2mp_io_d_out_14),
    .io_d_out_15(c2mp_io_d_out_15),
    .io_pool_v(c2mp_io_pool_v)
  );
  FC1 f1 (
    .clock(f1_clock),
    .reset(f1_reset),
    .io_d_in_0(f1_io_d_in_0),
    .io_d_in_1(f1_io_d_in_1),
    .io_d_in_2(f1_io_d_in_2),
    .io_d_in_3(f1_io_d_in_3),
    .io_d_in_4(f1_io_d_in_4),
    .io_d_in_5(f1_io_d_in_5),
    .io_d_in_6(f1_io_d_in_6),
    .io_d_in_7(f1_io_d_in_7),
    .io_d_in_8(f1_io_d_in_8),
    .io_d_in_9(f1_io_d_in_9),
    .io_d_in_10(f1_io_d_in_10),
    .io_d_in_11(f1_io_d_in_11),
    .io_d_in_12(f1_io_d_in_12),
    .io_d_in_13(f1_io_d_in_13),
    .io_d_in_14(f1_io_d_in_14),
    .io_d_in_15(f1_io_d_in_15),
    .io_wa_in(f1_io_wa_in),
    .io_wb_in(f1_io_wb_in),
    .io_bias(f1_io_bias),
    .io_rdy(f1_io_rdy),
    .io_done(f1_io_done),
    .io_d_out(f1_io_d_out),
    .io_v(f1_io_v)
  );
  FC2 f2 (
    .clock(f2_clock),
    .reset(f2_reset),
    .io_d_in(f2_io_d_in),
    .io_w_in(f2_io_w_in),
    .io_bias(f2_io_bias),
    .io_rdy(f2_io_rdy),
    .io_done(f2_io_done),
    .io_d_out(f2_io_d_out),
    .io_v(f2_io_v),
    .io_fc1_done(f2_io_fc1_done)
  );
  FC3 f3 (
    .clock(f3_clock),
    .reset(f3_reset),
    .io_d_in(f3_io_d_in),
    .io_w_in(f3_io_w_in),
    .io_bias(f3_io_bias),
    .io_rdy(f3_io_rdy),
    .io_done(f3_io_done),
    .io_d_out(f3_io_d_out),
    .io_v(f3_io_v),
    .io_fc2_done(f3_io_fc2_done)
  );
  assign _T = fc3_counter == 16'ha;
  assign _T_1 = fc3_counter + 16'h1;
  assign _GEN_0 = f3_io_v ? _T_1 : {{1'd0}, fc3_counter};
  assign _GEN_1 = _T ? 17'h0 : _GEN_0;
  assign io_v = t1_io_v;
  assign io_c3_v = delay_c3;
  assign io_pool_v = c2mp_io_pool_v;
  assign io_fc1_v = f1_io_v;
  assign io_fc1_fc_v = f1_io_v;
  assign io_fc2_v = f2_io_v;
  assign io_fc2_fc_v = f2_io_v;
  assign io_fc3_d_out = f3_io_d_out;
  assign io_fc3_v = f3_io_v;
  assign io_fc3_fc_v = f3_io_v;
  assign t1_clock = clock;
  assign t1_reset = reset;
  assign t1_io_d_in = io_d_in;
  assign t1_io_w_in_0 = io_w_in_0;
  assign t1_io_w_in_1 = io_w_in_1;
  assign t1_io_w_in_2 = io_w_in_2;
  assign t1_io_w_in_3 = io_w_in_3;
  assign t1_io_w_in_4 = io_w_in_4;
  assign t1_io_w_in_5 = io_w_in_5;
  assign t1_io_bias = io_bias;
  assign t1_io_rdy = io_rdy;
  assign t2_clock = clock;
  assign t2_reset = reset;
  assign t2_io_d_in_0 = t1_io_d_out_0;
  assign t2_io_d_in_1 = t1_io_d_out_1;
  assign t2_io_d_in_2 = t1_io_d_out_2;
  assign t2_io_d_in_3 = t1_io_d_out_3;
  assign t2_io_d_in_4 = t1_io_d_out_4;
  assign t2_io_d_in_5 = t1_io_d_out_5;
  assign t2_io_rdy = t1_io_pool_v;
  assign c2mp_clock = clock;
  assign c2mp_reset = reset;
  assign c2mp_io_d_in_0 = t2_io_d_out_0;
  assign c2mp_io_d_in_1 = t2_io_d_out_1;
  assign c2mp_io_d_in_2 = t2_io_d_out_2;
  assign c2mp_io_d_in_3 = t2_io_d_out_3;
  assign c2mp_io_d_in_4 = t2_io_d_out_4;
  assign c2mp_io_d_in_5 = t2_io_d_out_5;
  assign c2mp_io_d_in_6 = t2_io_d_out_6;
  assign c2mp_io_d_in_7 = t2_io_d_out_7;
  assign c2mp_io_d_in_8 = t2_io_d_out_8;
  assign c2mp_io_d_in_9 = t2_io_d_out_9;
  assign c2mp_io_d_in_10 = t2_io_d_out_10;
  assign c2mp_io_d_in_11 = t2_io_d_out_11;
  assign c2mp_io_d_in_12 = t2_io_d_out_12;
  assign c2mp_io_d_in_13 = t2_io_d_out_13;
  assign c2mp_io_d_in_14 = t2_io_d_out_14;
  assign c2mp_io_d_in_15 = t2_io_d_out_15;
  assign c2mp_io_rdy = delay_c3;
  assign f1_clock = clock;
  assign f1_reset = reset;
  assign f1_io_d_in_0 = c2mp_io_d_out_0;
  assign f1_io_d_in_1 = c2mp_io_d_out_1;
  assign f1_io_d_in_2 = c2mp_io_d_out_2;
  assign f1_io_d_in_3 = c2mp_io_d_out_3;
  assign f1_io_d_in_4 = c2mp_io_d_out_4;
  assign f1_io_d_in_5 = c2mp_io_d_out_5;
  assign f1_io_d_in_6 = c2mp_io_d_out_6;
  assign f1_io_d_in_7 = c2mp_io_d_out_7;
  assign f1_io_d_in_8 = c2mp_io_d_out_8;
  assign f1_io_d_in_9 = c2mp_io_d_out_9;
  assign f1_io_d_in_10 = c2mp_io_d_out_10;
  assign f1_io_d_in_11 = c2mp_io_d_out_11;
  assign f1_io_d_in_12 = c2mp_io_d_out_12;
  assign f1_io_d_in_13 = c2mp_io_d_out_13;
  assign f1_io_d_in_14 = c2mp_io_d_out_14;
  assign f1_io_d_in_15 = c2mp_io_d_out_15;
  assign f1_io_wa_in = io_fc1_wa_in;
  assign f1_io_wb_in = io_fc1_wb_in;
  assign f1_io_bias = io_fc1_bias;
  assign f1_io_rdy = c2mp_io_pool_v;
  assign f1_io_done = f2_io_fc1_done;
  assign f2_clock = clock;
  assign f2_reset = reset;
  assign f2_io_d_in = f1_io_d_out;
  assign f2_io_w_in = io_fc2_w_in;
  assign f2_io_bias = io_fc2_bias;
  assign f2_io_rdy = f1_io_v;
  assign f2_io_done = f3_io_fc2_done;
  assign f3_clock = clock;
  assign f3_reset = reset;
  assign f3_io_d_in = f2_io_d_out;
  assign f3_io_w_in = io_fc3_w_in;
  assign f3_io_bias = {{144'd0}, io_fc3_bias};
  assign f3_io_rdy = f2_io_v;
  assign f3_io_done = fc3_counter == 16'ha;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delay_c3 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  fc3_counter = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      delay_c3 <= 1'h0;
    end else begin
      delay_c3 <= t2_io_c3_v;
    end
    if (reset) begin
      fc3_counter <= 16'h0;
    end else begin
      fc3_counter <= _GEN_1[15:0];
    end
  end
endmodule
